%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20220919020035Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R 6 0 R]
/Count 2
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 7 0 R
>>
endobj
5 0 obj
<<
/Font 8 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 9 0 R
>>
endobj
7 0 obj
<<
/Length 1032
/Filter /FlateDecode
>>
stream
x��XɎ�6��+t�ASU܁ �mI���� s���)���I0 ����z��M#���h��$�yL�������ӧ߆��߿�.���c��1��Ç�����w�_�q��4�N�&�}�$!C�y
)љ�Cv�&�˯4a�1�# ��IqQ����@j`�,��/��-;�����4ҙ;�g��ɕ���@m�!l��_a��]݅ssn"+��dK��"����Ex���3X�����(��%�i�j6��+dC�Z�b��3�T���l � �3�S�g�@Ŷi���`N�~�#���lF��X� JMπ�p$m�{�\�1��Ԝ)
��C�xr!���.�mj�⡍R:wA07M�`4�g$�[4��Lf��0�F�f�Ʀ�ׂ��Z�4x#>�,1ogP�Yd��3���l���iI�_ٌ�a����(�[{�@fc��,�X��s����	o	��g�ū�>�%U�]��������]I�����އ{`�Wo9�5Vv��f�{*��q�.j=���&����~�֦�$B��j���H���B�FW5í�Z��Ф.2��.{�9�����:GW�.2�~q�,�B�׬;%1)W, �sV	5+�
vi�E�j�V>}g��]g��[�J� g0<�<��7����{�Hft�mOh�v.K�s Ɂ '��şZ�ӛv1S?b�m�Rޱ @C�`cg�K�V�/�z ����>kN䲫��%�zcӦ��Q�~�I��Rƚ��������
��j���x���9uC0���ꃅ�H?��y��]qY����HW$�*���� ��7S��:{���~��5G�=����Ѵ5Μu�g�ZR�\�'�r��/g��6᫶�
�#�h�˧��B�A�t'@���o����gf���
��X��׆f`Q@��*`c���G������]EL}�yE4S�h]��$Wlٺq���*�:>�!��������Z�$>�7���E9�ܷ+RM��u4_���bq���/7W
endstream
endobj
8 0 obj
<<
/F1 10 0 R
>>
endobj
9 0 obj
<<
/Length 378
/Filter /FlateDecode
>>
stream
x����j�0E{��ʼG��"���y@�@���GaSl��Y�m��ƺ̝+�2���3A�T�!�꘼߇���&}�h��6<L�Z.��rM�s��cBH�����v@$ �BEB��#���>�����8j�y��� ���ZU<��=��X��,y�`����ʉ�����#1-m�:�wF��6����#��EW��e�H���-�
�׌D�Ff�"Q�$�lsd��@T4�@8�*�e�(�������!��B���8"�,ሸwq$�DL�刨��ގ#¸�#B�ő�,�u9����ێ#캄#l�ő��J�r�%N��0��8�X�p����櫠:w	�P�֌	�8F���oѿ2-��ZUT[?�r�����]��
endstream
endobj
10 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 65
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600]
/FontDescriptor 11 0 R
/ToUnicode 12 0 R
>>
endobj
11 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 13 0 R
>>
endobj
12 0 obj
<<
/Length 505
/Filter /FlateDecode
>>
stream
x�]�͎�0��<�����k`F�"e���E�L���"5�Y���s��J]$�ח�'�����0�K�m�cX̹�9����s
�~Ȭ3]�.i����<�=>nK���Ze��x�����S���_�.��p1O?�Ǹ>ާ�W��a1E�^�.�c�������\w=�x�_�q˿����ӵ�J;v�65m����UQ��j�_ga���W��r:�?�9��XZn����X����r��d���k��y݂_���Wּ�7ʲ��	޲���Z�N֚=��ȶ {0��2�>���>�����OKy�_�?�>�����?2���
L�R�K�|,�k���G&��z:��8���ӿ��K��Y.�OG�
���^O��\.�{�_!G�R���п�>�w��Q#���PR��YR�o��7��ǹ����{�,�/��п���/q��L�L��w�,�~���,�������K�
����8��>�qu�u1}����q�.��� �
endstream
endobj
13 0 obj
<<
/Length 11059
/Filter /FlateDecode
/Length1 16648
>>
stream
x��zy|SU��9w���I�����7�^J-P(��6�)-BS���C�(��0
#��� )�P�*�#������2¸͌������9'ii����~�?�M�g}γ�g9I�e�iQ+b�T����q�\g¦�E!���sC�B����s<u���q�R�2w��z��x�!4Pl����y�0��:�1��w��������ީ�z'�������JB(�����4/�Y� u�ɷ�p(ԯ!�Y�����;����-��@}=B�2h��!���3,�
�J�������l��b�����s�kPrJj��!��Y�9�y��Æ�1b䝣F�)�Ƣ��/�=�#+���~7Y�b��/�Z����HY�!����2�z����]�(=�Z�~��C����D��Kh=:���h�{�,��-��?��_D��ux��{pfQ
����.�ڹ��2tBoa��3[���������c�Et/<��s;i`�A�1cP�[���5L4�kOB{�,t�F�A���vZ���¾=����H�}0^�6&��>4M�vb`����y�m�z�
{�f�8��z=
���Cux%ډ^��h;.��h��}�?�2������W�_��5�24y���37���A��I��07���!��G�Z�bg!C�@Ц%������9��-E��J�Y��S����h���U���5�[U9�b��ɓ&��N_r���h\�X�`��Qw�q��a��9�Y�i�)Ƀ\��8�Ѡ��h�*�B�9��(C��0�,=>W��W��!�5ef�<5a�'��ť�JJh��k�p
�|}�k����m�)���qE�p��E.�ϜR�E.��L�i�K���8�0�bE��ÞEm�5�#nרǹ��ՙ�]���J�4Ws;N�i�I+�� eY(-�Յ˧TٝNof����UD��8
2,�+(H����։��m�;hNM���U绻*��`n[�ֶ:lLv�/�"(��3\E��t�tj�:����a>��۾C@����-�h��l��b��S���{��mm��i�i�ut��q�W[�V��\�F�U ����u��g�7l�i�#�Q�=SK��)���L�Gl�A|\�;�Nc���ԍ�-���Iذ�CBs�n�R��h����ӽa���t��X+IOkOO��ȶ���-�%��s���­s@����a��v���dGd{�X�_�(��`��;�Li3Њ����H1��. C���k��Eq @F��GaZUX*���J��='f�j@`�ET��lWs��*�.A�����N�N[ƅQMmtV8���+����(���Ru��/���`ȽEd�mhYJq[U]}�Qc��}W/Vٝa�����^�v����T9�TW�U�V�J�̬�#�H���㒋o㪲G�����J����^h��W�(x��J��p�J�p�X��g4�,����H�P��Ӹ�h��q%v���23���%ajIO�)�P�~�+�M��qD��*���u5�a����F�C�e�yTV����0؄���S!�{��}����{�%�u���۔�Ҋ6�� ��aDTX��h���lh�^� [�n�vI"��a$�_�檨EG�=y����eB��tZaf���v^3�]�k*fV3@̷fZ�!3�j
�탠��N��2��4��H*�T�(�x�1	�V���Z�����){�0��`"m��B)t!	1��Ez����)#m���^툰LR�RRIZ&���c�tZ^�U��a-���v�5�6w��v�d��h�R�5�����YuX�`}�B��u�k a�[)눢,�6��x�fC6|q�ƀ�\c AV���a�������H�@���؆az+Ⱦ<��̪rN������`T�_fr+��d�@�@I�V@
�JO����g�&<b��mt�渍N#�4:W��J�2W�L��B5<	���i8�A�ѫ�l�1ʞ�N����|�Obr��v�����K�"~&�!�T`4�"i��qHg�1z�C���:K��h�qH�$�EB��K�k��eA�b��*3*H7"w\v�=��+pg�#(�&��&�)�`r��8Ed48E�"�2x�Ka��;���?�_2q�bŋɿ���s�^��|u�c��x�`�����=(�W��IH�bQ�d1	Z$��x��ܫ2��r/k�P\Azb�	&vh�k�`�� %n����W�߯_y}��7o޼s#�K�ǃ���x�k��?����?-����NE��@[j*(�Ñ�W*UI���.�̕{lz�A�w� s(��+(p�݄C����D����4Fp1��CSݱV��γ�F^�5�͘s�J��
O���IU3�LZ�rQ���c'2/?u瞮g؊ׇ�ȩ�]S7o��?te��_�� �6:,��
�r���!H2�qH�%[��^��U�g��c�yn�=�;�ʔ�΁�.[�$&�mv�K���#�A��\���~��en{�'^��z�C�����}�8wm\c5p������ӏ�~���d��;e�:id�>>��LM�=��kJ��5�����@������񼆍�OL��{ZW��GS�<��"@#ZUN`z6�(�R��Er�p�����ҁB�����Sz�&'�Ŗ�7��
$r�Ew�����ޅ߾4/��A}</}�������2�Ģ��ހ���ؼt���x6���`pZ�z�]�*�"���T�sN�ԩud/����P�K��T�l-P&H&�H�)��ړ�ĺ�Q�a���w�"�T�a�y`st�CG�wm :�g��|��7��a�BЋ�4�!�M*�S���h��T*ޠ�#�܋�*�}y���Od_���b��S��	y)Y����!�X9K1;!��=)�Ь��岻~u!��5�x��	"{|� .��Jf��!_S)yn�,^���Y`{�uԮ8n|��ŋ8]��Փ'��h7�u��4CƫT�U������j����=<
�j~�?�+,σ=媽�骪���kGЈ�}��?Q�luF��춮4fGW����̧d���Mr�ĕ"'��)�c�4��X��at������ro�Š�(��uV�(��\�p�z�p���G/��=�twx�Cc>Uል2t�p7��E0G�'43s_<��a����ܗ��}�ԙ�^�d��K�Gέ�]��\鑫�VƗN�w�9wf��ٱ�ї�I;l�ͷ?��}����<��`y��(��k?�*�FI�V���y�^���j��R�ǂJ�֨�(�/��~n�?��n+����������w6n��&m���3���`+<�o,(M�2���f�"��'ơro\��` `0��r�y���
X��:dϞ�G�}�J�J����[5������Ϭ��=�錋�^��x�9��<S�������3�?�S�	k�C�L>�?<�$.!��p�
�Z�`ɢ��Zm�:����54z�r�<z�wJ���Ɲ�Y��y�{�KiJ>���zv����d�y��ڶ���|#=�A'���?��`�a�� c��m�F-�|���bb��z��;*���s��Qs���7��7r	�啾G���������8A�jcWhr���Yk�0;#2�M��)���j����d�c��	p�j/g�9_�c#D
�!%���_>�܈���x\繫Kw������b���
V��ƷXMR�rЋ�ې����IY	�ZS$JH����8G'�����R�^����l��{>�,��[f�Dé�h�	�Od�:�M���o�_A�?^>�a��>�k���"������ix6�)?+?�b�ɟȟ�?b��?��� �и̅��;�0����K4(Y/�Z�ޡߩ?�����jV�g�ք�ת`UAo��U�(�w���d�w�Q6�7�jN=�0��ǝ��\�����~��X�S��7C�y��_N�Z�j��ֲՓ������u��a������G���gN��n������ M^�,J�����L�g��@��z,��6����-���Ĉ�n����#QK�V�j�eFoPA/P�����gԦ�OMJl��s"p���AÉ"�M�/>�+�>�}��]�B[V��({���)�;JAyh�4"Κ�N�I�������C��=�`�V'I�&'�F�#�5*؜S#�2�{�^{�I �-tg������CI`���AaM·$"���Z���Y���7�	����3�ۚWm�t���׶-ǜkǆ5۷=��f���O��򈕳��<gW��i�}/�8k;�.p_KS`�ܺd庖���7�G��`�$�E�%*,:ˀ���QM��	(�/�#�U?�����cpO$�f�V8��s�?�s}[kˆ�˕7?���m��t2\��/W�X��}�}���\�g��Ǩ<xe��P�deXV��t	�5H�T�J�|��N`W��e0���p�r����r���W����`�� u͍�(5�.����cF�b��c�,-�z�C��h9�lA�d=�����n-���|e�
;ٽ�t�0��Y��� �Y�zv��5�q]��>��߇�E���A`�2$%)��A���J�H5MƠWn�5�X�N'��I���ج`�㚂�����
~I����^IE}�ogް��Y8���ou�Jo~��n�� �_�}�_��雦>���ǵG,�z�O��v��z���Ɵ~��t��#xY@w���^XN䌇��ۀ撨��%����F�J� m��,�f-0�:�^���V��yk��{I�vnvz_
#�\���Q 9��R� ��pt/�|��%+�ႊ����ܗ{(����O>8��g~�b>񑌽�܍��u엿�1���{�w�[\��3/���jo��P)A����j���xA��W{��`���v�
�����N��t	bՋ��������v���O�Ķ?p��K�?~S��џ��v)��J$��8��l�����qlB<����ݝ�Vg,1+�6=�#�m^����n%XP�.6%�H�Ͷ�� ��e%Ǟ�ϛ&q�.�f'd�+[����Jy�m�w�o� ��h�z��O�El� �A��I���0�_F��,p�i����L#�9�Ѱ		6�.'��j��<�߂5���(X�MD,(Ʉb�)H؁�n�?�{��Ν��a����Ʋ�N�?LحY�����?�i*����u��_�&Ǐ��x���WXJ&lUbs�MZ�z�!��T$�(8�G���B���e7b��A%^���J�D��d��g�. �~� �Ϙf�nq0���þO�i?7o�ԛ[��7�bk������Hi@�0 �tzA�d��R,�j�6����d�o� Qv4�u�D!�-�.`Z$��y����K�=��,}6�a^�sB�_?����O�^�rc5�q̰�s��go��Ӈ���O�ǯ�|�=��1��r�����ũ�F� �-ƪD���i�1�D)�'17�s~�r�hR;�٥���FvMݱ4��	�<�k�g��a�@l�����77d���yJ��)�)�$�0�bm������8/o�o�����q�u�\é����œ�7j�g�ͬ���1D��}�{��� Z�J*�GF�y1�FL)P�;�<��s55}i�{��M��`�`�����=�#Cl�������+qF�JZ�`��)zE�	o���!IG�������� �?�?F�(��j���Hm�a�G!�`�,"�D^����tY�!�b���: `��"�TxWD>
w�xqW��ׯ�d���+7�[����|b�C�V/e�_�_u�4h���.�ޱw��u���O>�û�������Qj��bľf������s����iT,�e�=��l��3@�g#�¡X��P�0j8f���շ�����)���(	���hf���Rb��u�ӏ?����'b�Z�]7b��<�E7���'����@[�/��*KmC+�V��ʥ4�]�Tr�l�s6H}�Ɯ`N���͐�hd��
�[8pN�zE�CizD�Bx���Z�+��4�_ۼ����m���gL9������_y��e{�M����Βk�-K�K)���s(�ʑb9�l��5��fQ[�r/�0 D�����a�Q�x�{d�:vD�6~��9B��3�;���ve�F��Ű�j�j�11F�f5�ը}��� _Gdo�Y��쉮�tA����������w��8ԕ�-��4H�1oR�_(�`��6P7LJ4Z�h��f2VxMH�+�B*�*��ѣ��9)�>�e�#�)z@�]x�̭���ɍL�;�$��a�q�����9���,�
�"�s��d��cS������2�uB.�r{o�����A`��&�U�x6�0F��B���.�m��ʋr�;l8p��۲�4��ix�i����o<��}$�<��j)�Ĩ�V��T&��T\�M˘�j�d֛
L�I�U����jt$��wl��ʛn�`���x�Ɩ���z̾.?v�$���_������|�mz�)�z�/~�'�$t�Ğ=/i%��sC��/VR�Ĥ�Fx9%���� �4�Ms�2)���X������d\�Y=hT �ZK��%�
��*X�o�t��:6"R#�$@��d�t�}����+�����/�At.�ՃT!�0,�O��+����� g!
��ĥ:��$��ZO��aT��#衄�u� a�c(q궮�kOa���vh�����_ɫ��^㎤~${����}��4n!%
��
0T*�6�S*�@��� M5D}S�^u���A(9�{�.�£n�ƣ�S@��ow��b�y���`M�3�)�o��x��*��1K�o���������� F�$~Q~x/Vɧ#��7a�vͣ�L� 9E� �	�@ۀD-B�6�����g�������JB��k�=-qg����s�,=d%������/E�%��M������%�����y=�v�o?��B����_��ZZ�nYuQ*n�x�'�\���Su��8���i׶�����G��&W���M��� �2���t�'���Φ�,"g��t��IfD�3v���/��9�����	�-V����8�\�%����x?�,�!� ���kq��~����_XyZ~W~��'�����[p=����h���1֮��7�%ȏQ���,.|�.�n�5j��I�+;��I�1ƒ��jo\�T�T{5%ǀWd�=�]�nC��:�����HV'�hv�pb8��_��'�A�Uxf���>�+�˒?��~�<O�����ߺ>"��]��F���#J��*A�2�
���bU��Yq���D���/n^���§�Yu-��E��7�ٹ�#�C�ayvиx����I�c^;�U��+�
{��i����M����5��;A} X���iJ�����P�Ȧ���m6Y�7��m�
�Og6�H}��G�v��W��J�U�e����]��5��g����_�g4�O�Y==���rx�6B����T�
<���JN�E*Vఒ3�AA I�S����rS�_7S�'��'�sg�6y�Y|N�x�-bp��ft�[��Ct�{`��7�uA�R���X�x�aY�6F��0���l�2wl���%�n"��/�G>)��&�)�3��r����"&��ɳ�s]׻>$�e:��C� Ѳ�Wk4�K�ӫg�a��9�`�u�����n��:Ot������|Y.�t	����vIG�/�{�k�jp
�|���3}��&�m3����<�⋧:���X��w]�'~�`-~����2
���`�P�(Ja1�?;fq�M����ĺ�Դ�$jT�U����ӥ;9�`0D0����&n'w��XN2�J :����7c��8�?����?$�c)�<��k&O�;�~~s �9[�e���l�ؐz�����8Brp��� ��0�d�P � �6YK�ӟ��=�=bt���^�����ϼ�<��SO�{ozJ��l�wJb|�8�����B`[`�@7�@�
���V0x�<��d�<�w?%?&?�$����D�O�<rF@#�K4F��_��_��+(�t�֊���Q�1������셞��vߐgp �����v=��o�����b�,Z�'A�>�
բè�B��v�M�y}�N@y9ڀZ��oFO��0j��D/��Ú��>0vC�P�B��F�����5h2��zXe#l�A�<�~�Oq���g�<�1SȬa��u�������q-�~^͇���w�	�V�BP�*��LQ.Q�S%��Ta�9�u�0��ך�*�o5׵	�2��q�1E1�b��L�]���O�������a�a�a���{�!ʡB����ʀ��ݐ�c� 1қ��z�8���顆���-���Ώ�9�H��#z"Z��l��@�P{��Dث��
�@�#e5���Ѳ%2�����b�E�1(�UG�:���9����h�$P�H�A:�-�h(�-s0�-�(�{0Z��3ZV���kѲ���eJ��-����o�e�C���e-�[e��c�<ՂhY����\�8�1Ը�_'��B>�6м��qnCHL�,����ws���q���@�/�h�R��}X�8@��B���ڬ��9��Xqb�)0�?w�|_��`�����"f����:��$弬��,���ۆ6E�j����Z����[�s�!466��YYb�/�o
���:qZ�������~�X�o	�`p � x�[���k�%��z��Ê���_�����@S�/kf���M�qqCcm������ƹM�=g����>���)��.�i-�����i��5Š���>
B5�B���PKc�o��� ��0u�iqc������N�/ޗՃ0�+6.hn	,��fk[��&X�W��8�1�|-�Z`�6H���}M��[�~@v�]e�z����tt��_$"�R��$Xx~ p/!�>�hօ2��]h
�Ԁ諫ځa�څ���ס�|�-�k������P�ydv��ŋ�|Q�Ԃx� r�/���6��"i!P�/h"�[H�L��_&Nn�x 91: C�Q�ܬ������P0+�8?+�27{���F0�`~���Q��A��Z��h)�|2�ZE���ᝇrP.�"�F�>��8(��,��Q�Ԅ����?B˃��(%tv����Z�P��@o_�"�H�:o.8���ۂƢ ��CO�!�L��/�N�=���<�(>Y�$~n�/CmH"�q��,P� ��_���TnA���Z�J`W
:���$\�՚�i?��dX���R������.D ����<�uŠ���-+�;�^+*(v��i;�i_!ԃQ�"<#0R	4A;��b����@�>��:
�hXSt��9���s}Q�4Q�-�b�(��r=}�M��e�Z����߆�H��2��}���Zh����ݶ xYuNt?-�����~2+��I�^�H%ݟ7��j,Y��m�4��h&���O�$%��s`�|�n��'>*eT�!�}��T���iK&�Z��G9;lE��B�p����̧���n���Ѷ@/�ɨ�ѕ"ϧ6��^)�S͋p��B������	EWP����{D�0w!�bdgE�:�o��Q���m
EqY@wJ��f4��l��|��6��?��ݓ�9��z���r��.i��e�X�M��oa���#�
�Fe�r4G���x�wn����^�mTD���!�O��2��0�'�
e�X�^�L��\cSp�WQ%�}O�Ӑ9p%��ܐ�T�2x���h4�Q0~$��:y�㡇Zhl�p3�΂7*�y`j[�Ꮄ�¼h���i͆Vx#�5pCO��T8�F�8��h��8���c�� �{  
�]�@}�4�u�����x���q\��;6]�y��6pu�U��U��*v\���ʢK�%F}�����)������$��<���<�gX��cs����q����_`��a��8�qlAc�	�5K��l�����t��J4քm���@�Axb ˊ��f�c�T�v;���U���ϵ������V�����[+�bO���(Oq4��≜�'���'�q�q&�x�������Hq�9���<��/��<�c8�ţ�G[���r�G�G���W�8FJ�W�ho3�pg��0�}�� ��@� �y��L�����Ηp��1cc��aЁ�i�[��*����Ѽ�}rk��מG�6i8�jK�\T[uF�3[F9v�U�b4
t��ۃ���:��n�~��-'��Җ�i���ޣ<���W<~�q^�*֢ �J"�؆ǣݎ�q�f�؜��	l^��A���M,��sS\�Gܘ�����zC`����;�g�g����pk�
ʁ���ĚC���)H��gݪ��	�kV�v�~h��	ݎ�c�C�C9�9����J��A>P�&�p\e�;�R�f+�l�U�}��Vr�xhAr�=��,q���û�Lx��L�<f+�<4]y�>ʡg�1���;�xŦy:�ZJ�S�펫S��0Ҕ�;<Ҕ�4����|.�p�zJ��.��@��������\�0�����<k��+y�Jv���h�s8��j�
=��g�'��M���n�� ڮ�� #�w�0�;���i���aU��0^N� Oi�̰�&�*gΪj�x���P��p^EU�f��4\�Z�`�nC��`(Z��p�D���i�����{.L*8=
�-0j�����L$c��` k
�B�A~^0�,
�q�iAx�,	��	��{��zL�.����`�Y�^q�o4c
endstream
endobj
xref
0 14
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000392 00000 n
0000000115 00000 n
0000000549 00000 n
0000000604 00000 n
0000000761 00000 n
0000001868 00000 n
0000001900 00000 n
0000002352 00000 n
0000002779 00000 n
0000002979 00000 n
0000003559 00000 n
trailer
<<
/Size 14
/Root 1 0 R
/Info 4 0 R
/ID [<BB7AD869AB7F21C58E803ACF99B92F21> <BB7AD869AB7F21C58E803ACF99B92F21>]
>>
startxref
14710
%%EOF
