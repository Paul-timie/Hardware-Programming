%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20221103023811Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R 6 0 R 7 0 R]
/Count 3
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 8 0 R
>>
endobj
5 0 obj
<<
/Font 9 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 10 0 R
>>
endobj
7 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 11 0 R
>>
endobj
8 0 obj
<<
/Length 1113
/Filter /FlateDecode
>>
stream
x��XM�6�������KU%X�{����VʡRs���v��M�H	~��<WS����U�v�VQ�"U1M�߾\>�������K���n��M�����U����9�����_/���)k��ɘ�N�w�5.��%�9.�8_s����pq�΀��Y�7�T�F� 5�Ý��A�K�S�=�o����uxq�b%QW]�p���W�0W�1L��p��=�9O�t3KVp�����*��3�f���졄��t+��1�D�����}[�A�� [ ������(Ց�9��}�A ��椉f���}����CȪ���j��p��f�6����J�C�C��?���F75y�vS���bEܳ�`Pnܣ�xNX�Ĕ�벥�(̇Z�~K���KԢ��Lj���ԋEp�~2g���J&��ݛW<(��oB�F�<..��qO���<� z��L�!a�r\-^�%a�N���1i�|V	�4��)@���K���w;+� Y�(�.���Jnb{�,*���9i,c��E�C�EV�0�`Uоß�xA� A9ތ|;��������EՄr�z]��q�s7�g�{�q)O�?78��z�FC�/N�%)�Ϛ�'bi�� $�Tg�8;ʠ����L�(��;o��!m����ĕG`���x�!��%��'���yk܌,��D��
|�|��rqzѯ���ם�/�&�ht�c�Z
k���:)k��px���,��DP{8�v"$� �;�_���\u���,��qb����Z0{�j2q�ACP���ԧ�h=D�V��G*"�>�o��Xn\3MS�K�\Qn�a�>#�g���~���}��J{��#����O>a՘vcZ�Q�,����;i��>k#l#ei#��Jb����K7U��� )���{����c��h���tr��V�&�G?���|,
�9`/�Il��zRa�-Ǘ|��%�k�#�iװ�Ll��N��ho[(�y�;,\g�N]�0l<�WP�&IO�0r�G�h�^je�vR���aND������7�<БM[��84|�o���y�	y&\%Ғ�����j�l#�ͼ�Դ�ܺW$&�\��a�ɔ���?��E�
endstream
endobj
9 0 obj
<<
/F1 12 0 R
>>
endobj
10 0 obj
<<
/Length 684
/Filter /FlateDecode
>>
stream
x��XɊ�@��+t�A��7/�}���9d.��T[c�c��4�	��zկ_U��vz�a �}DJ�>����G��S�8?��ӯn�Br�(�?}�?O�#���_�(A�=��#�E�+Ы#q����O݃	�a��p��a���E�O"M0��n�j����I�ƅ0��-��ԃ$(Xhd�	�_�)�tM���&l��S���А���`�D$�$�	��< G��
�2�$&�k�d�<H[
�Вފ�s;k����	!�r�Ի����W2�w�z^��� <K���0�ǉ!�+O�hiy~��YBA=�"�BR��k��ЎHr6��I�������3H&эB�l�w/o�[�]�������<BY����K2h^֠��8G��6��S���8�Vo�@[���Esu�g*!��VH �iwW2��3+���]�/&�r�Vs���(٭�
5Q�-���(�ib�[
q^������I�0��]iɳ������}��`a��}!`���z}�n�m� �je��_v������#L 
3*%�!����YAL8j.��L��pPbIᥪ�YDE/���(��jH��G`�?��j@��x���i�vpiz��v���(:j<ʩ.��@�	-\�2I�ߵ�����x�~;�`Ԧ�E�s-p��F��j���Z��
endstream
endobj
11 0 obj
<<
/Length 256
/Filter /FlateDecode
>>
stream
x����J1E���Z���*�ꀸ�Lg?��� ����-i�=�!�A�s����>	�(3��LZ������c}a�����R��d_hy���Ġ��	H��l�������ŝ�N>_b�J��	�9#�}�!����n��l����W�]��>]q�'�6Z�Ru�)M��i���$����;��;��h=��8�8һ]��l�5�j�E���_ 2�af�V�`�l��y���H-�ѐ���D߿��P
endstream
endobj
12 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 69
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600]
/FontDescriptor 13 0 R
/ToUnicode 14 0 R
>>
endobj
13 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 15 0 R
>>
endobj
14 0 obj
<<
/Length 523
/Filter /FlateDecode
>>
stream
x�]�͎�0�=O�r��}L�)�L�,��f� ��!��}}�q[��D�6�/�l{��~�~�c{�Kz�n���>�>=�K?$Ʀ]�.�H��k3%Y{|�=�q�N����m��ӦO�K�}�;?��%}��=���}�>��K�'u�v����Lߚ��t��������+xL>�zlHi��ߦ��s3\|���:]��u��k�CN����C�	�ynwuȖ9G�N���r�\0k}���������5+�f� �r�y��
yǬ�o�Z��<6d�3;d��f�C����/p�E�_p_C�� �/0���I�����c�wX��~��_�o�/�![��,�e�L����_�c鯴��k���觍����_�`�/t,���O���F��D�����K���,я{I�?�%яuI|�[�������_�?B��я�K|4�o5�_���
}�-�B�U[���9�-���Ը�����
��E?z���
�+�"l3|�lߴ��sغ���=������d'���o0E
endstream
endobj
15 0 obj
<<
/Length 11269
/Filter /FlateDecode
/Length1 16980
>>
stream
x��{y|SU��9w���IW�B��Pz)m,P�P
�mhSZ��6Q
�@Y�QADDIQ�����0��������,l����}�sr[Z�����>�~I�g?��>�y�s�p˂ ңV�"�v��y�iE��aK�°X��y }!����9�8r�5��M�^�3oq�A��u�����l���~�(��]0Ɛ(�޹_��C~@���j�^-�o@~ü`�����G(w����ۼ���%A^l���'-��7C�(UFhD�on	4_��}�a|~	�a�����3,�*�F����&��j�;b����%;EW���Դ�22��sr��=���m���G�U(�.S\��?��g���~��Q���pÑ-B���u]ꪎ�������T�����kh?څކ�CJ�j� z����:��G��1��G���Ga��4�U����^D��=0�0ޫ�.܆YT��h9ꀹ˹v�M�]ćЛX����V�a+���o��Q���#p�N
�oѣ�(��<Ö�5����߄�'�=x&�4��@�j�3V*;�B�AjA�~ōv���A��Ft���(Շ���u�j^D�i����>��9ƨ;G��w|�P^�v��r��m�%�m���Z0���
��ߡ&T�f#/��FS��,2�H������i��kʇ��L��A����F��+���s�����7�bT-,�������e�ƏA.^ܐt����ʩS&�O�8�l����wxK����
G�q��a�R����������2���匳�MFC�N�Q��c�2��)��)���w����Y�bI\CqVf��[�b\�������F����߫�&"A��[ZJіROKlG�d
�9W�;���U�^_�����4=���T�����=(U�Z�$�]��VR4�v�v�{L@���ڵ:H� Iw7���Q�&�����Rǐia�%��H�䪒�D�˗�96bp�*4��DTtH����֊�'��u���}���gU��C�6���mUĜ�.�\�e�<�t�D2Ȩ���3��8§��b����|�o�_)RL�#��0c"xJ��|��u[��-z�j��]��ݢ��֮׷5� ܨ�
���zembĻ�1�4��>e��)�#��3�"L�Wl�C	��]�%��=m��S5X @��"0���l�DZ'WE�"��xI9�SCjNv��+IMkwMO�7�v|EU[�K[�.���#��A��ƸM��.w��,��Ѷ"P5��Q�� ����ti3ь���r"L�j����0��]R��-l��D �4#*S�"R1$$�±������5SfFr����������Ɗ*�E������Z�W$���X�VS%���\uy�.�_�!��Ǝ1 e�%mUu�gMb�]�X��H>��]���^H��ᣲ2�j|�{��U�)�D+�p\J�-ø��À F�)j��Id}����p��R�p� pZJ�h�X�Qwk #2P,	+�H�Ϡ<�1�ݣ	$�)Mt�\�OV&բ21�PPK���LA��sL)-"X������� F��*�6EY�b��jj�\/� &���3��H�n���ɖ�R=��ZlS��W����ʀ(AD���̉��v��M��T���%�(s�p2�{l]���jm����%d.��O-���V��ƫ'�KxuŌ��&��VO�:�`fLM��} �UaӠ�)%�$#�i
dԴ}�Q	�VZ�����������0��`�e��D�t"	1P�Ek������e���~��L��Z�Hz&�IlǤ���>����8'�C�)����k��h�Vh!E)\]ys��U/�t�w���|@\��ٰ���uDP���j|DِX8�ݣ�M�Q@���h݁���]D�Iya�\ �*Q��нx_�DfV�@%ńӉm�˄S>0*m�����e��/g�@�Bɒ^@*�jO��s9��<l��c���z�.3�2����r�2W:-�|�F5<��>�4�8����+��1ʙ�A���.;�����v�"�=]�����@��l2	*U��c��d`������j��l���+H��ra�.�������i��0Ì<q9�wͺ�Г�� 1��k�X��&�'��X�%"��%ZU��ݟ�ß�����|H�I��������z���0����5����Ṹ�i��G��L�h�MD:��%�E�#��k��>�����X���
3z!�M�g&dX�������� ����/�����v�5�oߴi��L2L}�����_���������@���:�;�H�ii �Ng�Q��$k��9+W�Kp�&�ѩ�ȡ0?������z��������2Gi1�̓�<�v�(��w�F�4Z�X�FK��	�	L���UӭLz�ra�޼�E�����Χ؊�-˭�US7wƁ�w��{;׃��^��sE\9 �F�I���@qҠ)��r����W��c <A���E2���?��P�Mf�����H���J�;,���o���7^Y�ඇ~�%L��3�'e���yj���/>���>z�		P+�v5���:ix�1>��NK�#��gI��X�I��`�����]񼎍�OJr���Lzw��G�}<�֓E�(F�@N =��(��������v��?5�m �L-0�-��Q�Y\�6GJ�(<�,����*��n� �n_��.�֥���c�x�ۧu��f˔������fSc����Y<w����Uf<��v9�|�p�S ���)S�.�2k�C9R,a��@�m��@�l��� �"D�JO2�Bņ�k-����By�m����#�W�޹���9lҹW��́��@.�Јv��h���d�i�f�à��&���>�U(ٜ�Xȃ�E����B�=�;����O͞�6�":��3U���m��t�*a��<.���M���[���o��1�B�a�dX�5�����o�	f�G���BX��7/^��G��܉]D������ti�� V�U!Vë�}N>�g�p+��e�A�<�r�<����A����!K�Aâ���(f��R����tfGg����'d�梍r�̍G.���Rǲ���������K4�R�}�6�!�ܧ5ؑ��'r��q�|0���[��n�
�;4��\@E8j���2��a��~�F�03g�٤�=w���x�[GN���,V�=/|�����%�y���^��my�����7���,lk�X��Oި���[_|ž���'�o;X^}DY#`��V�b�ɩ��a��x�`�i+|:��e���cA�Y��c��fT�����V�3�Ko��ʯ���~{Æl��O�����
/�%�IRfB1�*�jUŰ�Iq���5�`?0��l��pU`Z,Zbrf�����|��Rk64�&���Up1��us�'<�y��K�O/~+�<��gJ��?�oB�ҕ8[�;����q�����R"��"v�׎J6� [��k�Z�)>�Ig �[t�����4�O~,go�{ꭗ�OW��5+��٭�o_�9浲wjۚ���������
s�A���5���;�P�,6@��+��� k��s�H�V���~/������������8A�zCgxRY�5�k�0;�<�M������NΟ���T�&��}����j4��S`M���s����c񘓟\]���w��|X�Η�G䗱�׿�Z��-0�\��@v����X�2�ѤB>���
 �8����!�*��v+6�����%��5>�"_|xV~�a;'�����^������Ϣ$I���l<(@aa�Uł]la�x��_��H}�R�;	�0��$��RvB���h���1����I�xg<c����h�!�F��C>6�V��pl��-�B]�n��[u//(���w�]���~�|d��gټk���"������x�!?-?��c���_�?aÓ?���8� ړ@��%���T6��_rL�٬��*��z�݊o����(<t��u���MP��eߔ���Z[��tخ��ѕ_m{g���`��O7,;6=x�������d$�ս{��}���I�+��A���aY�\k��!�Z���g����m�X��pYrڱ��t��W:�:�`���m6js`͉(壹Ұ8{�6-&��?&&K���<���53F��2&>N�M�2(�KIa�f'A���7�ч���8��%�8��F5�zA6`EPJ�&{2�选�޾����|���}ͫ�g\sv^[�ퟭZvߚ���s�X�z��G7o�K:���+�۹��g��=��Ego���ii
.�[�]��e��6���a��4np�j�6� ���cca��bC>���4�44^5v-k4�v;Ȁ]�jB�fU���������u63@����Pj�a����9
s��מ�mƁ!O����~���ڵl�֭�e�&2'�g�Uk�'Fp�3森s�S�:��ڍK�6
>�Y��]� Â}x��C@+�*��j�^������X-��"�A>��Y��)�)�`�����*��u�n��`#��m�<����߹C_���~@^����U�pڇ�_����@�x�+�JBqj��c0X�؄xN�3Z;�NJz��ԪV;��A!��Ce�gO��0bAź��4+�*�#���g����ܳ�Y�Dn�����̣f�VսS)�ÿ��^�������f���׫Q�y �M*�(R	N+�/������;XG?�����0��rb���K]�y*��m�^9�lD0i���6�F��~'Nf�{�?�vZ�߆���><y?a���E�Wܹ��Sp���uN���4)~��`��gZf+�mD�Ù>q���1�XJUq�t:=��e�K0n�pZ`T�j\�x���UHn}b;�3�Q��^	�w�h��c����rc_r}ælA�Am]_s�8 �.���!��(��vR��>���& �lwl�z���9)���8iPl�uhQO&j]ٻ�v/>s�^�tü,���?/z��u�[u����1C��ކ��n�7����>��_���;��Q�����8��i�v;8uvG�]��?�`s��(�;�2���X�����zz�g��Sv,��bB7^��*ͳ��2��/P��t'y��L�QX��C)�=%5-5���fG�#6-6�����{;X��?�q�asL�6�8�7�anĆ�,�US}yC���z� ��]+���%�#�W}�3�+P��<��Ojj���Fu�,�GJp�l0LL|��><�{o�ģ�9�
�l ��@ۉ@p?�3�/�����.}nP򑜆�y�"{��T����Q?��fi7P߁�l+�Y;JF�R�.�@��51�s���u�kB��jO�B=��>�ͭ�g�&��s�#.B�J�x0u��O�.��kr:ށ�ٴ��#�m���gN>�����K_~���%{�-��wϔk��-���S�����\)�c�V�Vg��6�]e,�q*B<"�}O!�Z�T���x�}���m�;��0|�������v�t�0g	̹
�W�K	`�F�e-��ic���!6@�gD�{ǹt^�p��$�e~��<�֛�Ӱ�4��Tб`!�F��[M�N+�I�L��#��ƛ���V�}jV�P7�'��.6P��|N5�v�^��#�_N�W0{R��A~�y���SM�2_��r��G����l1�jd�HIf(�^��s�ς��rl�����Mf磖� ��J �_xwҞ�����ɍ����Nz����+����0=���� %� ��6dKLj�bd5Yk���V�I��a�%&&�Z�qq&�dcp���6�X��I��&1��NF�M�V��jB=[���@�>.Z��k���t�Ժ��͛=o��x̢S���BL26���f6����ss��k~��bT���R�Tɢc��(4�l��8�Ue;�_��n0���tnߎd,b	ހ��(_�g�c�:��a{��r��Qa�W��;d(H��d�i,9�3��|ɍ%�^l��"k�+6�Z*@11�׳��e9��3�\&Y��Rh	ZNX�Zx=k� �7S���q��ޖ��M�oD&�wN�@j���G������ګ�ƛ~�ߓ��qg
;_�K^���	�ϳ��˃Z�Y5=��`�b%-KLe��N������ ��Q�H�˗I9�(#�Z9�1�I��F�� f�,��K1�U*T�S�|o��u���	�HD����̞�;O��q�d˓�_�%;�y)�r��H��1@��������v�	�3�K� �in@������{\��׮�`T̋��7�;���|l��m�3��/�;r�C�q�e��;��<{��ǟ���z�������U}�FéUj���ꐮ����W��*
�`�#�3�P�q�4!���cC�x\#?�Z���\)��O��'�5<�c���>#������c:	��R��Q~h�ȧ��t�f�vΥk�x7@\���I����/I�P��粲����x��ׯ_<�j�}�P.0��Z{�O��!9����1p����f{���ݖ��&s\���O��qG�"�w>3z�C�O��2�/>��y,n���W3��]R]��[:���)�,m�V��6*�l�«["���G#��wΈ)Md=��7e�9%�9O4�7���"9a�|��^�� {��E==��3=p�j�>�Z�}d�?sfV�L�!bM�k�������O�Rp��������'z�O>(o��x:��}F���;/��ʗp\T��Q�%���0�&�x�֮��$$�;����c̥q�վ�8F�����tj��Q(S��2z[l�W�QB�K �	�c2�Qn�W�Р�<#�|�{��ŏf���=�Cx���ɇo���/��q�.�k�Z�Ĥ3�|sr� �Z,�6 ��g�#���hY���h!�Q�ͬ^�Q������X���Y}�	Iq�r�N�*TD�XQ���>�$c�7���@�K���;:��#�?8n���X��P�><߉��v��~}f��w6��h��������L��+���6!��<6��B>5o�;�9�����N09� ��z�k���٥�+k�`�������7�z|ʯ��u��7�c:��o L��5�ɬ� ��jR������9�4�!f�����_޸��O<��8����w1f��x���=�^2���A�R6F��xX-V�VūX�A������h�-�=�ct<l��G�m��!�s���=�'�kc�H��Z�C�ZI�;x	�_g7K���#�f�Ҭ�^_!ƪa�D�Ϭ��;�tO�?��57�K�Q=-����1 ��G�$�Xi83:���<�Rs�=Ұ�՜EJ_D���6�o,肆�韇�����'��6y�9��<�[��Υ�����7�י�t��`��������5�
s�t�3,��Ǩ��@D��{#O����v����{��ko��r�8:-��|L.f2�<?�y��}�O��>�a'��Z��caGP�Z�%*ǝ�^M�,��Tr�8��y���'�������|Y.�t	�
!���<����A�FJ��4��`�H���������F������F�\����f��G�GW��2��y,~7[�go��9�s̹��<5�@JP�\,hu˱�����A�[w�a�"�)����m3��s[�9�yw��v͍?����ݘ�Z����؟Ìo�b61i��]��ɓ���=u��݌M��|ǥ��p�����\F����c�a�S���E�A����q�2��df����ˠ0�⦳���>M���*����|F.�m�vr9>��$���|����f̕íG�{�]���Q���=���W���F?��j�m�B��;��=?��؛��y#�����9�~�h���I=�M���Y�]9�HP�1�8�/��2�$��T`�� �D #s<�>da����g������'�G�G�s&�#sPADQ9T�G]�»Tr���y����>`ԟuQI�o*�����	F{�	v>t�a�Ѓ4��ӹn=*���ca��u���g�8t�(�6�
���ٌ���;?�yh��@���d�˟�cT�A�0�<���q��[^����k�q���e�!_^���;�㱝�y��ߞ=���?��|����\��5����(������ġ���ߊ��. �� Ŀx�qpݛ���:G|L;;���rI����=BON~oQ� �nC�ٮG�r" 8z�kM�iU�q���3�[��,y����]����l=?��<G¾��{�d��^̝C��DH݃V�Z�j����h#|Bߢ�ނZ�R�	=	%��r�����X�u���QT�0J���a�7`�3�M������;�]xX�͠u,h��	2VG�> ����'<�1SĬf"�5�������s-��K��k�����)�I5[��TU�'�o�?ӈ�4�K�A���7���%�Gu��E�4���+1���1{z�DC��c�q���x�x�4�TlZiz���Y0W�W�_T�"���7�&���D�=ʚ���67��:�c����J/
(i%�yJ��6+i�cJZ���JZ���v%�F6��Ѵ@D�i-����%1'{�"��DIǠV��(�-$�s�`}J�d0V�4��[I�h0���9hP�<J�T��w*i�ƽ���(�?��5(�����2_��)i�M�?JZ��Ԙ�t�����h��ōsÍKub�?�k�͋[�4���ځb~n^�xG08g^@li��Í��l�[��S`�R8S�T�]�8;m+N6��,��o�4�Z�,��d�ZB$������YyK�Ɛ��-���|��b��/bK`Nc(h���&�2�"[,��Ma��T'N��8����6@k-a?4��ιZCu��d�Pv�����	�p8
6�C0P6&� ���54�6���!�.j��ճ�}{�P��45 �[K��%jhl�#��M!1hi�W���0Y��@����?o�b`��f�:���1�@�oiJ'��� �`����-���ЬPmK �������5�a���`�kC@Cl�7e�,h	6���w��l�E!�-�h�@�.DXRK��`�y���dI�� �.ܐՋ��`S�E]� �.�O�X����׶��y�?��e7����sr-Z��W�S�Ɇ�s~�.��9�����2^�@���d����e�f��ĉJ�L�[<��) ���p(;�8/;�2'g���F0ύ`���P��C��Z���b�H�(Q:��g>�Eyp��h��y�_Dc ����O��&��Ø��h����PQJ{gBj,���ʠ�l��=��&�g����<�mA�Q�����Q\�<�/�N�5���|�(�ٰI�\�_�F)�aZC��O)�ʂ�q�"�P���&@sutT2v%�����iO�B���D[M��'���п��e-��Bt� �<��-��:گ{m!�����y����-�sN��$�uE�)�bF�X@9���E@������::��&��l�9����~�7M�sJ*����=D�m�9DH��EJ-A��*D���� ���P�mk�||+�60��:[ѧET;z�OzE1��E����}��JP�"�dV2n]�MD�(��z�J��S�=��y�t5P9�S.��)�ݨ�)�$s7Ӓ,p�9��d��`+�~v�(z���pf�7�k�&Jm-� MZ�Sf��x�Iw�p��J^�::Z����bVfR����{T�w�bT��r�7��ߠү�ڦ�B�|�)T��pp/s�:�ͦ��[j��Vh����G�j��֒�Z��e�h�ѿ�4��`�ʨ�hV�ǫ '�2ѝ[�g̗w�*����0�'D�̦k���`���/M?�L��|F��
��'�J<EyN�S�9q%<��<�T�2x���h$��~8<o�<y���Z�ht6� ��\�P�A�8Lm+�1\��<��F�c���9P
O$½.���.Ҕg¨�gI�/�.g�h3.��5
��H�B~�4�u���ӝ�zӝ��r~�-pn�����+l��ƫ̉�x�U�Z}5x�E��K�������/S�_9��՗�N㗸��{��ϱ��������ąw/���J<C��q�c؆Fa�k��#���#?��l�'�h�;�"r�ay�aYvT��06Kl��S�I��I�'��D>ጟ���g���7��ɞx�^��l>����Og���g�ǜǘ�c�ǂ�;�?�B�S���(�h�h��ɛפ�@����i=9µ�f�/�t�%��H�K���M&9y/��,<��z!�s��^`r`v>�O�o?3:Q>6�:�Mp�p��
�d��;jv4�`ߚ���7ՙ�M�� /mu$y	-�����-#��Fkp	2v����)���Xb�Ӹ���[XiK�<��ő7��kܜ��p��W7��W��^�Gק:��r�߄s7a禜MLpӲM�h�(nd��qI^qC�f������l�:l\�\����֙�^�	��U�P.\l�I�;+z���Tn�y׮Hu�7¹z�H窕#���r�|�V�+sW���e+��B����?A�&�p\e�'�R�a+�l�U�u��Vr�ziBrZ��w�(u���s΄�xZ�-�<f+�|$]}8q����8�*pJ��M�v`��N)Ot^��5��&��&��{�-���p���s���Yށ��x�c,V
�p���ޫ^�Ջc��ґo�4cc�)�Xɀ�aЯ��:��Xh�6.3rFc�q�1h�h<o�2�
�쪑"0x��oj�Z��1�C�5e|DS>3�WGR*�]�<#"����3��1��{h�zT�o|$��*R��7>R	�$Z!a���@E�P8^��`%B�0<i����2�?�dpF()%�r���
uw$m!�`>�:�3B�!x@/2)��aD����=%�tW(��ٻ�����C�]�(����'���\B8
endstream
endobj
xref
0 16
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000398 00000 n
0000000115 00000 n
0000000555 00000 n
0000000610 00000 n
0000000768 00000 n
0000000926 00000 n
0000002114 00000 n
0000002146 00000 n
0000002905 00000 n
0000003236 00000 n
0000003679 00000 n
0000003879 00000 n
0000004477 00000 n
trailer
<<
/Size 16
/Root 1 0 R
/Info 4 0 R
/ID [<B3127F0E3187F00D137E2D64C7202E93> <B3127F0E3187F00D137E2D64C7202E93>]
>>
startxref
15838
%%EOF
