%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20220929002115Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R 6 0 R]
/Count 2
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 7 0 R
>>
endobj
5 0 obj
<<
/Font 8 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 9 0 R
>>
endobj
7 0 obj
<<
/Length 1099
/Filter /FlateDecode
>>
stream
x��Xˮ�6��+���Iɒ������� ����������X�|g� !��c���C꺖�/�4�q���tDm��������~j>�o`}��2�.�kS�k���{��B����/�~������|�|ʚD��2&��]p��.����b�o9+f����p������笋˛����Z#9\����I�S�ή�O������k�'�E��������+Lg��ǰ�.�	ל��y�i�Ւ'q�4���zf7��+,�7�w�`xx"�+*�1�F��sq����H�b��\3�8�J1r4�Մ�ϻB=PB �掫��N�$i�qY�N�VX�8oviS�]�0�g�QN@3��S�}ި�.��a���R7���5e'�#>[�NHK��¥��̇V��ֺ�Q��wZ�O���%�~2g	�_%�|J�&���f�2M����((�W�$-��I�(h�r��"�W�J ���Ϲ�&�<�Ig�� �@� ����K�v��|�R�5��>>���L+�`g���Ni,cp���!`Ѣ�7e��
�����f:Ǜ���c�Qr 9`�"4���CD�t�߆5<k�N��yr����]t%�5�o��`I��>���X$�Ag�:me
�Z�dL��(��o��I]��_�F &���*�'1��E���t����nF�<j"a��!_�\�N,S9;ſ���&$�����OH�`]e������,�DЙ�����&���ڟ��K���]���e�t��hE`�v���(Al�<���^��y�������9g���X���#{�q����h33��%F_U	��Ζ����T�k1򌛲*��X���%��V��Z���\z�ln�(,���Q��yh��A%u5�~MEV���a�f����hS���.W+"q�>��1�Xm�_?�L{?͢����#8�{�h�� ���DFaw�b�����F����=p"0�6�wK��O_[��$uF�����<��Q�2{}z�+ _<0���	��u�B�@��0 [� r�@q�����6RX��wg@�t~8ᐍ�.A�h�Vj'��$��'�b({��j?6G_|j����
endstream
endobj
8 0 obj
<<
/F1 10 0 R
>>
endobj
9 0 obj
<<
/Length 336
/Filter /FlateDecode
>>
stream
x����j�0E��
��P�cA)4���}@�f���$n��R� �-�֜�{ǰdޛ7nM$�I�H�����ʼo��?7��	ѶF8�d�s]�L�t��pآ��& # �nÝ�<��/M��(k�8P��0�j���TS5��:}�q�C���4�%�1S���
���2eͦ�"�㘥�&�b��/�+k���k��Η?
�_e����� �V���
/S��>�{b�����TOȪ�`?%�:O*XU�B���Zu\U�9�.+g��2��z�,Z5��j�S���.���t�Y�����r�h���A�k��~d�3=���
endstream
endobj
10 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 65
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600]
/FontDescriptor 11 0 R
/ToUnicode 12 0 R
>>
endobj
11 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 13 0 R
>>
endobj
12 0 obj
<<
/Length 502
/Filter /FlateDecode
>>
stream
x�]�M��0���>n�Ğ|�J(�C?T�? $�F*I_����33~<0I���0k�m���_�y��ߦ��ys�aL�3�Эq��ݵ��4���_�y�l��{xv[��y����JүK�a����1���y��~\M�Ե��9����_ګO5��Ї���x)�>�7Nז*�����v~iǋO6YV��~_'~��{VL9����Bm�2��;r�\��r�d�/�+���o�/�w�+c^�[eق�X� 7���;�ƿ�5f�:.���9���2�>���:������u�/8��_p_K�������_h��>X�W�K�w��_s�?j:��8��o��%�\�r����U	��~��88�8�ѿ���5�����/��5��9z��/o�������?ǽ$��>�s�Yb�Q_�_�'�u����G�]�_)Ge�;x
�E�/����5s�������c���3���/KE~�AL�0���y����ߗ��
endstream
endobj
13 0 obj
<<
/Length 11013
/Filter /FlateDecode
/Length1 16576
>>
stream
x��zy|SU��9w���I����hiKC�"�Kic�,�Rh@hC��2��&� #��*�(� ���(CQ����8���3�:¸͌������9'��e����}�|7����9�y��$��%A�G-�ER��@��cEp�A[j�FĺF���1��5-X���;�!�mEH��E��l���B�"���j�z�0��d��_;:P����#w�ي5P��k�j�sIe�5�.���X�����XL]2���-o
�#3P���mHSs���o����+�Ç\z(
�ΰ/���Ng0�����OHLr&�Kq�����i������34�;,/����n=fl�4�~�g�3�|1��j��sq��-C��"�u]쪊��Y���X�c��+� ڍނ��J�ztzu�~
�Fϡ��ځ6�a��q���������:އB�.�ֽཌ��V̢jA�Q;�]Ƶq�˓�|��5�n��<
8<�>���}�o B��/�y�;H�5z�����b� 찚�ͯ��S�^<�k ,����Jc'�u�n(-��ï�цt]� ����݉��J��mb]����Qڶ�{���mbN0���Ѓ��ZT�W�]h�\/�D;p1.F[����V���d������7�MB���?SS��2�H������i�? ה���L��A���*W��0��9���#��h9�Vs�����J��U�Ǐ@.^�!��9���3ʧO+�:e�҉Jn��/'�3��Q#G�����5$s`zZ� O�+�f6q:�F�x�e0����8ʦ�f_�S�	���ꋆd{|�Q1 F�ťyJJh�'��h��������e�)���&q4M���ѳE�ϞV	�ME��D˓i�K��8���0�bE��������Հ#n�i�{��C2Q�VE��=Mmx�XL���QmRǑea�Ł�hٴ��"����9!j��.4���
�*
Rl ��b[fG��v�_��������������3��<E�A+>O�������h�Z:�g�қK�(�j��"؎��ž-�EH5}�H1ʌ���nr9}@��V�G��V�ڻZ�{D���M�om*r��J ����gԷ�5U��Q~e��Q�9�Q&�'�������3��?u# (�v2lh��|�D[�U��"��<�����&=�=�
�����3���--�l�r�j=�@��h�|����1S����i��ő�~:V�&�6�Q>��zO �!SZM�b�.�����q��8Ş�j廴> �@蒌� ̨�JEP�
Ǌ�r�aF��PD���4Em������+�eZ�6>��k�Y��b�WbqkuQ�3��8�v�o&:_��!����� eiŭ��uQW����N�t���8��T�D�B��;�p���̨,-��N�]9BA$�A�q�ŷ��T:c`@ ��T�X�8Y?4A�胂�p4<��T5�& 8m%�[8Z��N�=Ј��E�8R��'�4���@� g|���wǮ!�t���0CM�Z��f
:� ��Kh�ez����=�bT*�${#�TV�Ai��jF�Z/b����+��Q_��7q���zO���	��b��SZ�J�{�0�ED��f'�D�=`{E�4U��6I"�\?� �L�m��W������ҹ��eA��tF�L0m�m�~Z��חϮ<n��o���#f�W��@_�q�meH+i$�T��PQ����B-����^ӎmSw�aT����L����Bb����Hݣ9hS��Zh��!���%����L�lä���1���8;�`�t�܎[�4�36�FH1�W�\�bv�z��*$�KB=0�J�XKe�����O�9�5��Q�l�D}T�	Fu�B�^@�b�iW��b��-���(&0��*)&�v��.N������ȭ����Y�
�Hz�XĪ5<	³�f�5[�ȑf��;4�kv�Y�ٽ�eV�0���ia�6��)�=��	�$Jz�;F/��1�({n24��x
���۽�D�wv]�����$�T	H��O@��1j\&�7ت�f��CB� 	,ʄ�BT8/\=+[��XQA�y���ͽ������0��k�Z��&�77x<������,����Q�E�{G�zD>"� �$��U�R�๧�������7ⅸ�i����y�L6�p��MA:�J6��GJH���k/�@	%d�� 61����aa��y�v�P�&\���u����Wxl�֭[wmfR`�sx 6�x�(%������?�#�r��ka�tT,�w���P�\)F�Z��8��Y�2��h5�.d��^��P��X(q���1\��to��;{s�m�u3֡㤩��G����YVf`�biݾ��
'3�?~w���'��W�ʩ�[]�p���wf��}�:7A��^�gq�\P̃FH�R̀qҠ�vg��l|�N�]�� ��P���2����ǡ ��İ�K�B���*x�ps<���o��Ҋ{��]���+���o�����<{ ���$4T�?��Տ>��ͷIJ�Z��끾�!���F1&&Y��题dds�ZN�[,�dcb(�\�ĮD^�&&&';���&���ϣi~�W��&@cR�'=��(��������v��?-�c �L�3�ϣ�Q�[܄6Gj�X<�l����.��v� �k[��n��Ņ����Yx�[�w�O���'��,��TM����>����m��gT���䬲i��O:��L�^Kt���D�sʖ�	cP��m���d�����!�UzR�xo>��!�r׋�H��ះ0���wtG�&"#|�ȩg_~�3�.�x�f�#%�Ec`Z�Y�՚��FÛ�Fė��3�P ��71�����y��{�#~8<����5uC�E܁�sT�p�Iy���<K�NX�z(��y���F�r��'	��Ux|�{�.Y��|M��sx#�;�Y�QkŮ�n|�8C��5�'��h�u>��:4K��5�j�*���xu���g�|��?̟�U.����rU~�t5U~d�#hd̾ݔ�,��ʽ���9���Y�b�x�<�qٻ���h�\ɥp��2=M��Xv���F�2�r�:���2��d�,�kv�*�\�p�z.�pB��G��ݖdwx
�9��p�Ɓ	�?��a��~�Ac1�`ߙ�v�w|�}��7��q��g��j�9����>�»(P��'W��N,��o{m�B̂[sb]C e�>���7?��}�տ�:��pY�1e�@� ��FK.�^���y�Q�-����6"��f��(��͘>5�y��<���^yc0~F~��[�7ofS6���[�~�>�JBS����U�ժ�c��	�̟��5���LZ��N�"0--��s���mo�R�Rk6<�&E-f;��fp��Hz"��S�.\�ZN]��gJ��~����4l�:�?��%��?�K�<~��v4H�p�vG��je���&�Q �ܢ�G�~��{�_`��񜽩��7_t&>7P��V�WU_�>j��e�c^��NMkSSC��⠓]W���f��`l6�#ެ��PC?XL̲�Hb�*\Q֧X�֘���le���Qw�\VX���g��an�I�;#S'� �m̮��P�(Fjd&���i ��X��*p����Y~�W�A��kJ��f�=��57��x����{>x���G�|�|L~��y��%)h%��T�mH|�D3���D�%%$�3&`c�+��K����D����h�a�F���~6�V�O:z��Zh8�M�����,RAf��?|�͵˨�K�6�y���w��&W^`����w�<�ų��gp�v!�#�3�lx��^� ��yP�4B%�,��x�DR�bد7]�]���+�.��e�F�nO
��*V�7�ZT�JE��͞�w}��Bf���_-é��������X���]{����?�|-������ݫ�<�hˤuS�S�3�;�Q���Ũ�����'O?�a��⻩6Þ�`X�,��#�69�MQPЋ���7�ټ#7޵��c��g4�#�J�$�pC��f��K��3��a�Y����g�M�����u�X<|,�����&�X�o��][[�7ŵ�.����_mg���Ò�ټ�Ĭ�]���|���w��1�!�����kʔ�˪t�#��Ԫ�_-0�O]&��=&��7DN?��ם.v�Rge�e�bx҃ ��@����h�4.} �nf���?` ���t��b��`�X��u���v�T$�VCWUl�(�y3"Q���T�= I�bh� wn~ް,���,���)�+����P�K�q��9;u�gn�~�������.<���c���3��0�x����w���}�!á�^~vY4�3��s1�*�!�	V��fS��$5r��~���4��N'g�'��p_�����r�Ɍ>�W�W���+{�X���$h�J�~�㿾3��}�l�pOA4�uw��o��g���|���}�|"k8���Y�/��@�oZ�{>)]��	�Z�@���� ��.}�>���+�� ����yA|�Z��w�a(�5���������'䭲_��
6�+n��̎�,�U4α�aR���� ��ƛ���Zm��Y�BE����#)e�d�\N5��1�@�j�_��v
������;���ض_���)���&w^z���jX��-�HB	j��g0XؤDN�3Zۻ:$��\bU�F�@���/�1{��wo�XP�6-�
Hy���N��ϲ�k��X�p�/�g'e�+[�����
y"�Mַ�n��wd�F�Տ/�lȳ [ �JCS��*�e��U������"ܤ�$F�&%9L������,o����� �f$�A��dabA!���-�PNa��x�?�wY����7O��t���=���}[~ǲ��L�y�^��5s�s���qC�?s�*[���K��S���xv0�:Ii*��N���bm�x����j�D���X�xɂ�Ν[@}�OBgL39/�-���t��d9�-<8��6����k�jBE�v}�%�w@f6J�/�C�Q0zX����:��MB���c,���Bt��Sn��C�-�D�E[1�d�ݳ��x��2̋�AN��벵m\�Ⱥ��o��X4�ɟ9;~�u�1��}�?|��7�^� �H�ΥpB�&�i��!�;��jd��\
�cH(H1�	�/���G�*��ا�y��9}���n&|�P,�j��v��=���Ow��z�	�ħ(�����������wħǧ��q����aV>�?�	��Lo<�o�l��������CVMե͑X,w��	(���l�#�@^9�hPaF�T��:�l5. �RD��\�w%W�g ��A��u���`#��m�<��X�o�m�N}�v��!|���/��e�h��_���м�k�g��/�7�pǡ�["ę6S��Y���ϝ-@�����@����s��{��lF�</��qs���^���G�߷}�r�����e{N�>?wI�����3�O���ߦ<a��Pݱ�T&�9�pVp(I]�ΚdM��[���Xht���*f��i�9��6�[�lK���0��V�'ʵȗ���N|u��g�ɗ�o?�W�9�H��~�|�-0[�W�M����b�\-�n�K��qr> ���)�c�V�Vg��6�]e,�s*"�TL��R��M�D�s��9~T�6|�����y�m�g�{;��	`�bXs葖x�2��hYF��u�X!�"ȣ���KA�3����09`~��<�m�7�c�iP)�}�R�5*;K�Yl���˗��6P���;,�r�e~q5�4*G}s��|�
�ŴWI٢��N�;�ѻ[Z������_~?ɼ��}����e���#��|,	�K)qbm�ٜ�MV��&k����b�
��0љRb�&$� �t'�R�Rm� K�P@usoFZU7W�	��E�!��Gk0s�7�;L-K�x��_/�l>����v!&p���s��蓳���J|<I�kJ�,*�9��9"���+�]�������a��본�;wX�=q��X&WJd�3Z���[na9ex��qG|�p���7e�i,��fⱧ��+f���v��<��a�����4X�g�r.ޡg,`��Z��R`	YNY�Xx=D����T+c�ϑLKn�y:2Ob�bv� ���+�C�O�O�q��_�����Wqǘ��W��W_|�LR�s��s��r�NϤpX�xI˒#�Mc'P�*={n�!ab	���b=�0F�J��B+��ƽ�rLIa�w*��8O^��$��5>�*_X���=���S"���\�L����C�IR6&�#�Z9�2⩸
�F��f�,��J0�U*T�W�|�p��|��H	���xv����y�)�nn�ly��3����۰.�1�H)Y �S��h�q�Z��V�tU�N�z�PQ����������o�ƣ�7`�������Q����GX�r.�#%1�8^����v�Q�;�`78����>����cu'/�����t���Z��΅��S��C���&J���_��d���Od�j�~����KB��k�ɰ���!6�<"K�HŤg��bC�nKa�S8�^��y����чw==n��EO>0}�7�}p>�D��_�_��Y^�aEUQ:nnץ�^���W9�c\X�8���ۢ����K��O��鍰���]��w���K�F�����,���@�y�WW�l�%��$�%�\�d�'ڂ؛�
I�y'��K�����	�\���g-vr�c��,�x��ʯ�Xk��P�'�w�♉-D�	�&=;���}���#�:��է�州x�m�~�����Yx������yA�Z�y��-���$�_7�;M�Nk��n������Rb��$!�ʟ����qU~�N�1��3���(���&~=U�!J~�"ޓD��É�&�5���������$�(z(K����1��<S>:�o7�u~2X�e��^���|g��kNI Z��H�A_e��f�1Z�fc5d�zlf�z��u�<����P8��=�	CHÜ�Ӭ]Eb V��o>�(c�U\P~0��=������x_���ڎO~ c?���+忺�_]�Su靭��/+�ՙ}���a?���Q�d�F؈�jR���&���g���NA쎶�1�߸�ѩ%�?��$�J�����o:�k�����Js�3`2�R���a����2?�X<��Hb���:�T��|v�y�X�"���_K��r,�~�P|�=xc{ps�كq�y}V�\�f�O;��N��RF��xX9V���V%��I���S%&Bl�����1:�(���e���M�_z�K�#{�P�=l:�{�V�=��$���2P`<�ed���;2םn]��1^^3�z{C�WS=)?vw>�'�jX�2�jf"SE� x�vZ�ܬ�49xu5ϩԜ:N�4��a5gт� ��>?��'tACR�z�:<��<|Vn�7��˓ϲE�\�Y���|�y����?�_tӑ_��V�9�E:������TZsj���~����9�\b�<�,��{�S�+��]r��8>-��^|B.b2�<?�y��}�gBly7�d"�Q��q,x���E�S9z��3���I#Ǹý `�';����Ɏ�E�$]��_��ӌ�]�(������%��uZ-�`*�|���3��X�&&�배K���xc߾7:^����˷_�'~�a=~�W�I�v�87�; *u�$r���Rc�q_ ��U+H{��̠�$�������8k�k�=�~v�v6s�Y��q�!���h����,�"��3��8�Xj���������$��,�p$��9�W�&̕��G�{���ـ3�`"�E�M0��~�Vn�&�mۨ��߱��?ҳ�x�U��tɯJ|�A�������n��H��M�g���P�"�ڐ@mn.��V����<B��@��B����yg	N��s��|�dbЖ!���9�#�_FOF"��0�8����DH�2���q�������v�׳�<��=��O�t_H���X����[�>���h��;�T�^@-pB��m����kt�+�&Ԍ��'��-����Yx����l�쁜�-(� ���A$�6��X�:�u��v�f�����3qP=������@c���ǭ�2�(s��cw��s�\3w����!�A/�>UP�W��NP�TP_�$hj5��ڴS�k�����
�����������o�e��͏���a�a���\c�1j<o2�
MkL;MgL
������Fw@��5�Ho
n����bd�Vf�PP)��.R��Y��y��Q���R�*��)e5�����d 1���LV�:��t���>��X)ǡ<V��(�- �s�d�J�P�X�AΣ�Y4���9T�<J��U��w)e�ƽ���h X)kP2�'��e��Q�:4B��JY��И�rZ�Y��h��OE"+��bm kBM˛�Gā5��ܜ�9��ЂEAq|��)��4����o�+N%�H�8��&kR��`l�89��\�dQ�y\�&�Xl�����:3�&�ܬ��,���[�6�ŀi��!���"!64�#�fhlh+�ʳĲ@$���⌞�S��j���&�	��P��\���!\�PCVg��ߋ��Ҡ89�á��@��Ƈ��������zqY ,���{�r��,z�����R ��5뚃����b8����:��D��#�5�E���7�����e�z�~s`:%��@V76@�: �ذ��9��":$\�6�z�����E�Uh� ـv5aJ���hR��9�dg�>��@@/F�ph��`��nkÄ%���E0	^
��l�.�h�F��».���!1P[{��j�,&�ZG���4���iQ P���#��Q��˖-�
(���d���,o
*,i&P/�2�H���2�l�|�$qj��ȉʀL�[<�fU� 264E�Y�EY���S}�Pj 3� &�N�"� �P�ׄ���'��UD�u�s�8�[D�è�/��"�f�E�
7�Q8���Gh�P��`QBggBi̯�`�|��WD��;D�- ǳz��8�9A詥3D4��3iO��=0ʁO���̟�� �DJ��!X.����B�&�"�R���'Hk�*�]#��2:�P!BWk��f�ĊSa�:�_Cy�=���&���r�Bυ@�f�A-�׽�0�����i�(��-�kN���}�P+��ь�XB9��� �v=-(Mk)"a���� s�Ϯ%*s
o)�*�.UV#T���0]�����)��"u�`!R�(b|_�:���g��m��F�U�+���jg}��ɬM��{��?�t_��$�N�X�*��L�t��C(��~�KR
P�3�ucx�S9	P.�G(��T�UvI�n�-Ch�Lu>�Pv؊I?	1F��RJ8������b[K�B=�&�)+�v��ڤ_�p��J^���ڐ�@�:J���j�bT��c��K(c���ȿQ.@�R�5Q�QpYL5���a�e6`G>YT{�O��=Y
�����^M�������ŀ�$�4��ߒ^��͉r�F���hR�ǧPN�ѝ[��PXo�-��Ic�#�0�e���
+L�����=h��k\.�\k2��ӕ�L<ِW�����N�o�?����=Ə��mP'�<<�H����Ð	n��Y��E%8Lm<1ܱ֡0/Z���p�Z���H�g5ܐ��S�%�:�QE;rdye���\M�̸ �{,  
�]���>VZP�:�e]_�������sm������l�ʖ+̩+x��Ru%t�E�����������\_~>����).���g��\�O�������y����wϟ;�J�����	lCc�ֵJ�1lŹ1��d��h�; #r�a{��a[vT7����f���r�\!~\�q��я9���=��U�z��U���^ï����Nb�d�Ɏ�l�ɖ�����}��D����N�������������v��j��n�3�Ⱳc-ǢǸ��ѣ�������8)�@��%�5�D����l�����C�CLǡ�1�2����;����F���O�"�,��$�q���M;��Ms�ʗ���.mg �u$�.�Gfߓ�F�v���b4d�v������Z�#�.�q��m���Ҷ~C}�6�z���p���z��ü�%�G!��D�Mi�˻\�✭ص5{+ںj+�����[X��ᖄd��9g33uSզ�&6g#6ntm���JMV��$�"�9p�]Xw$^�'��d�mX��z`�h��uc\���Z;�˵�~l�O�/�>6�^�j��h��0�'��wN�H�&T��l� ����*��w�Ǫ#�4-H.k�o������9�ok����l�˂���:G��,>�q<������v��R��2��ʴ�i�4-o�O��:��n>7	O��s��J\e��)��� ��o�����]�1->���\{�+L��
4�~%;k].c��ʸ����ƩƐq��˨*��+F6��H����v��mFyFFi��kziTS6'��GS��S�6;*�����s*�0���&Tد4�[^���/��BA"�(���9P�?	G�d�.��(##�7���QF��Ig�#���3��XB��p�D2
��a��0)������Ȣ0G��G�� i^8���<��1\zp��a�^�^	�//'�b
endstream
endobj
xref
0 14
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000392 00000 n
0000000115 00000 n
0000000549 00000 n
0000000604 00000 n
0000000761 00000 n
0000001935 00000 n
0000001967 00000 n
0000002377 00000 n
0000002804 00000 n
0000003004 00000 n
0000003581 00000 n
trailer
<<
/Size 14
/Root 1 0 R
/Info 4 0 R
/ID [<D17F251C85982D53F3D96F1561E60CE3> <D17F251C85982D53F3D96F1561E60CE3>]
>>
startxref
14686
%%EOF
