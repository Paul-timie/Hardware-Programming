%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20220919020037Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R]
/Count 1
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 6 0 R
>>
endobj
5 0 obj
<<
/Font 7 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Length 895
/Filter /FlateDecode
>>
stream
x��Wˊ�0��+��½ɒ�����}@�Φ��s�d�Ċ�a(ۑ�s����s��𻣎z���}
܅T���_>t���?����>vA�>u���Ǖ;������?>�~���j�~��$����@�"%I�0�z��L�~��c��T]����w�X!50�*��'���ʎ=���l����p���SSt�����~���3���&�����&r��*Œ+8H¬qطR���Il�8Z�cv�:.�SS	��������ǭ�EW��.Z2\f:�f�큊��
�ZP��\���� $k��S,�f�k܅#�������(��X%Eh3?�'Rݨ榡�ڱD��R� �VM����dB��s�2� '�u���|�UaG��a��K�3���O2/6�����>Z&�oM�+g��@�2��1�+�-i���r0�*�YIYE�fF(8a��y��]�����J d �=����i�m��n��Ŭ�/�%4c�pa�l*��N�4�9��3/B-^M�0�S0�'���e��7#_P�G�!���h��\c�m�xV��4��=Jur����]蔶�Zyc'X�B�לOG�13�4e��Y&�ZYi�E��c>[sY��C�P��[��Yf`����k��D�Єz9�|��d)�%F[����%���i��2��<p.�N+ ��Q;&Y�K��"K��UҦ�Ik�Ե#�)�㦝�˂�!��d�Y���䷊����س�,�-Vw
@�۸�����:���&���t�'fP��r 7�2c��(@D��O`��|�57���h=�\j��5���z���x���M`�u���T���d�w9�:������{��m�8����`�+���/^�k
endstream
endobj
7 0 obj
<<
/F1 8 0 R
>>
endobj
8 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 61
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600]
/FontDescriptor 9 0 R
/ToUnicode 10 0 R
>>
endobj
9 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 11 0 R
>>
endobj
10 0 obj
<<
/Length 485
/Filter /FlateDecode
>>
stream
x�]�M��0���>n�Ğ$�J(�ġ*�C#�$2�����y�V�xl��G�|{��aɿ��;�Ŝ���6�C���_�1���C���~w�v��{|�=��i�����춄�y�������a/�������<��W?.�Ț����|n�/����|���<�cʿ����ӵ�J7��6���x�ٺ(���̏�guJ9���m��6���5�� �r)�R�ރ+����+�_q߂_���WƼ�7ʲ��~�2~ޑ5���1{�q�mA.��/��/��Ա�w��xZ�������/���O�J�'����^Y����M����qG�zN�5��5�k�t�/u?��.�_sS��[G�
���_iL��:�w�t�/����7Gyӿ��пB?%��.B�R���A����>�kݧ�J�?�(��(��)'x
�E����+�`N�����!���a֙�4��;��4#K?����&
endstream
endobj
11 0 obj
<<
/Length 10743
/Filter /FlateDecode
/Length1 16176
>>
stream
x��zy|SU��9w���I�����7�M����
�Ҁ؆6�eJS���Rpʪ"��*. J�:E��q�u\f�gt�q��EG��>�sr[Z���|���כ��{�{����o?i�mq�Q;b�T�(��}����SaKݒ����y�|!�ن��:|�e�����_м���/�MGH_��X�Կ�ZqBY�`��а�{� ��>�qQd٭6�
�?@���P]@�#A9{�/
,k]�5�P'�bK`Q00}�p�r�-o�#�P����m���-�zq�w�P!~�a�����3,�*�F����&��j�;���ɃR\�{�gHjZz��a�Y�9�y���#F�=憱����
�Η";���n�����'���=5��<[����
u��<z�G{ЛP�[�Z��@��^?�N���Ft�D����8��g%-mC5�yu�
�eh/�{'���w`բZ��`�
��{M.G��!�֠�p&�h؎>������&�=�~��p�I�o�}�x��<Ζ����Z��_�����x.�4�	�@Pj0W;�E�Aiq�~��N���G[��&t+��f*݇���u�n�E/ж�c�}l+s�Qw?���T�֣z��FOɍ�.���R�U���h_�LE������~�ZP9��|���M��S�x5���
2p����)v.2uiZ��\+W�;F��?��_C�Q���kD6��T�ޗW�?�xpCҍs����fUΜQ1}���)�'���+-�X<A*?n�cF�9�0?/7';+#=-u�g�ە`3���8�V�V	<�2e�Q\[eSE�/�)�ʲ��҄ƒ�R��6*�(<�4OYm��b�M�G�_smT�7�{S��)���M�X4�,���K<b�3�ʛJ<~1z����2�F+qPq�a��P+�F}K;Jk�Fܩ�N�Lj��P�VE����N�1��Q:��A�8�,�4P��Q]Z�t���Y��O	�B�QabTE���h�ؙu�cc�	ͯ���{�7WG� ��`K;:�F͙ѡ�����'�΃�,OIi4��:ef�:S�-��|��#v|�`;����!��"�(31�gV�����;:|��Q���i��M��N�����F�0EWϋ�Q�F�Tۈ�����fN�Zg̭�2�>�1 -�W�q�r��}�T��n� 8���M`��%��P��Ϩ��E4�yI���(SKzN��ثHO{oO��Z�vJeuG�K�T�)�7���A��xLQ��N���bG���"P5��I��i ��? ��0ъ����H3[�����S�)�U��4&�" ]��Y�Q�
R@�Xig^.��ÚJ(3���֨�S��]BViSe5���&FQm�2*�[J�J,�-��@��̨>��=g;����`��%�e�D���Ҏ������Yz� V;�Q��{��~"v��гN*~*+���Tz�̘S=J!$�A��RK���S�MU���j����E4�>(x���=�JU�e�i+��b5v�޷���P�4X��G�&�8M,�M U�gb���w�>�Yt���0BM@-��3j�ωe��`�@�^��=~O��*���<e��«Yj�����{+̨/���荴�W-��{Ro�ء�L�� �{�	P>)��K��Nj�B{���&Pi����D��q��3���SY=����v�
��M�Sfgg�i+���u3:%��rN��|�fUb03����9�����4h+CZI#���Bf�	5}�yDB���r����0�m��6�꺘X�)�P]HB�p���m�Ա�v�F?��@&iyI-i$=�8;1i:-/B����9=���N5�6w��N�䌽�oH1
�U][�jN�sz��*&��F`6��R���JcG��(r k�G�g<��3�Q�'X�y�I{i/���]"����+��H��j7���t��a�@8���a�"�[^5s�J��R��Ukx���=m��ѣ�^�7?�kv�Y�ٽ�eV�0���ma�6��i�]���I��bw�^��b�Q�L:I~.t��4&��g��o�9�-�� 
JEf�IP��^��&cԸ4Lo����f��<AX$T{��pV�Z�� h4l�_cEE�f�Mȭ�eޭE��L�yd]��� 6Y�#F�3n�MnѪ�����t4�w���C��L�\�T�o<�8�O�$_Z�y#^�+�N�s­w�d�k��I�4�C�(C�Y=PB��X�טX{��u I(�(�����zfB����,�m ��t��������_^��έ[���̤��g�l��8Q�J��O����}�G"������T�H�4N�r��jM�&c���r�$��j�]��

���^/A���Z(8�yns���<<�o����G|�A[c݌5�4}����n�V=��d���4<�?�x*��C�����[��Uy�j��9���\���Sݛ �F�ɳ�b��QҠ3P��4hH��Y�7ہ^��qW�9�����~$S݃�=��&F�@8��e�W���A��\����x��w���^��~�K������#8o]BS �٧�|�ɇo�ER��]�F��^�mLL����E1����[2f�-}�11�x&�RbO"�c���d��S���?ϫ�d �1)P�@�%;��;���"�`�]�NK�@ �
M�#�~T�7a�͑Z0��*[�&�Kn��+:�<��q~adI��h^���a���6�ؒ�������Ժ|��x��pgxV�y�SΩ�!���L�9�n��z��ρL%P�O�4�l�m6&p&&HEE�	��ғ��{GP�a��+w?/�T�a����~��^�ٽ���5z��^�΅��A.�ӌv��h�Ak2�Z��a�hx�ֈ�
?r�
D6�� b18���c/vď���!��r�oȳ��N`�\�P<�<�\��[+,Y���v�q6���\y��1�{�5�>Z�=L���C��Q��ι��s�,���bW�@��ܹs8S��5�;���Q�u>��:4[�k4��jU���������#܊�~�?ë\,σ=�j���jj���gG��}�&?�Y����QvGw�����|�.y�C�wMs���K� 7��)�c���x��ev��;���
��dȪ�kv����\�pA� L8��և��ײ��L=4R��80!�G��h������Y�ԩ�.�7���?��ï����lV�=-|��~����@�j�\ݱ:q�|ëbܚ�)[�#�_}�/�w^���3;V�V�X!�ՠ84Vr��z����:m�_�԰-�q,�4kW<F�@n���,<��^;����0���
���77o�̦l~�ĉؚw������P�.e% '��VU�LN@������dҲ�3�%�i� h�uȝ7�o��J����k�Z�vV����G6.ؙ�pֹ���?�;���z�.�)K��������+��i؂u�%*�I��|�y���v4T�p�vG��jef��&�Q X��q��O��ҽ�/0ނx��Z���;��P��w�46�ۭ߼$s���o�u��6��!:��5�#?�!9A���7���;���,6@�^�+��� k��s�H�V����G努�=��{��G��q����������s�ocv�x�(��R�Ff���?����'�j����|5��)���Ll칠|�܌G�Ix≏/-􃷙�����/���c�?�|��� ������h������Ģ��A�lLp%0q	�1ѕ�����1�רX{��&^��I�Aﯙ]�z�	7��~�E*�,7��o��|��x��G����=�������g坸�����1�	<�=H�H�L���G�k�^D�2��F�a�E�hH�Q��F�˸�x�x��c������Ia�]�j��VU��Q�����nc�3W`&�o$��2�
z��^��;��"��ˏ�.������a2^���ŕ?㿼�g՚�����Nc��O�k7�tFq��s����K�9��-Ko�2�{�m`Q�����x6DQQ?�ǃ�hc]}�Ɵ�I���6��� ?�����z�a�&���N����Tl
q�Ԥ��i0'�),2��o��T��=۰j�8p/�=-�mMݕ�{��P��;Q*@��	�lmz\�}p\\�`O����Y˘��6uX갰?5�5�]a�Y����ч���ٻX$HAl��F�0'�U
���=_�h�k�~�ۧ=�ֺ.�֝�O5w������U���X�9ϮM�v����xE��{q�v��l��=�����>�����Эm-�r�����n� xo�������J�jHV��A)qqf���'���x�«�"���#���H*��fX�o�����m��l_���w���ͼ�x�_6�::;���[��w"�b�ޝ��r�0Еr�AY��aY��%��!�Z���`;I��"��d��7�����}��b�p/vWw_�*&���Z��(-�.�����F�a��c�,=�F�K���9�l:A�d=������Xlw!��]����ۘ�~wT�*��e\�h#�������)�v���*V4\J�#����xXJ^P��5~5+X�6�\ֵP�@��d�N5��1�Y��{�ǧ.b��������l��t�|釯���#خ�����	�Lr8JP����8����&%r:����sB��eV��ad$0*(�B0���>�y-0-���i�V �ku�ap$�>��\{�?a���pĞ��u�l����������9���_�6=��М����^�ف'A/�@���I�T��
6%"���g���1�Ԥ�$F�&%9L���X��i�D, �m��9z��JqMB��D��4CMs������{����0?(����������-[�]��K�2>tp��Mӟ��'N������W��&�[�peL[��b�a�u*��T�#�N��!Lڈ�
�� m�;�x�7�����̛7����gL�1/���t�`��	c���yu_ze��5l-A�A=_r�`��]������`��!V���
�Nmb� H�7�%��cN�Д��M��th��{ �X��x���G��u�[�X>�</���.�羍kX��٦�'�7�߁�b�7���͟���/���ۀ�����|'$h��f��G�#ήFƟχ�9F�Bӛԙ��w������l��ǹ1�3w-��a�W���D��:O1�?�`��f�{2A�b����Դ��t�������Bv"N�7�:���g��8�>z�����͗͜r7v�w�ê���9���0�8j�ʥ\L�X���F<�`�_�p�zK��e�*��X���4�]Y��I��oǫ���7go��ɖ��?�\����i1��Yx�d�`�s���!����κ d)��H'�v��X�/@����/�aT̳��7�[�����|`�];�.g˟�_v�5�G��.��	7��}��ɏ>��[�aC�uFA|����8��Նl��V+FV����jm���
��#љRf�&$� �w�w�V���X���&����n��htkB}��lb~�%Z��˿=�|�Ծ�����M�f󱸥�/��1)��>��0����>9�p���7~L���w;�o;JAR��iP�9du:9��.QgM�&���VȎ,4
v����?s\�my�Y�*��4<&A<� �|񲜁w᯷�|�|qǎ3�Y3E�b��������zd��D�!�ٯ�ʵ��e����#�dĆ�x��ZmZ�Mgwشv���ϩL��l1�0P2������<G^аM_�[^���)y���;�s{#`�RXs-躖x=���hYF��u�X%�����l`Q�����A���������z�pO:����
�/a^�y�by6[{3��FH�f(�^��s�߂��
?��HN����9	�>�)
cFIPْ��Lߛ����������/��d�8�����2U���P�4ɢc ���#�ǖ~�ˀ��mg��\���]���۵���*�U
�DV�������e�.
V���#~�H@����$�\�Yx�I��ꊛ^y`{��<��p�T���4X�g�r.ޡg,L��-E���咅׳�y3��X|0��d���\;�y!1�!�J�}Y���q��?.�����]�k���A�������8���4{��<����s#�	�/iYr��{X�4vJ����C�?�p�(?�P�4Lǰ�C<QS0g4�0���u�9j<ܰз),�{z�^��!3�ɡ�u���1�8mG����c��wݻ��;�;��;�5|�O/q/� ����{��4-% '*0�>�S���,��j�;����F1hʁ9By�)���^=��ʯ����]\��q�� kQ���$������ܮ�j~�\��G���9@�|�V7 N�{��'c�nW�a�w/�{����,4Y����A�z��<��3X��&���A�9VS㗄
��ڗ�zs�C��yD�vA��=����v[
��q��?�#'I�޿��	�.yd��a�~��٬�	[o��(���tÊ��t���6nH]�xe��z��<���e�3/m��[����/Z<�cg��~z�����s�e�4,�B/�11LIS����?������x�#�d ��t#�ڙ�)9C$Y�����f��l ���������Ʌ#^c��k8�Z�'H�̙	x-3�g�5����\���~��\����������>���'���<� Qx\��ػ�����!�A���3�D�a�x���i�Z�M�S���g.K���'$0ju\�_�Ssx3F�La x2�����*�%?OA"�#���~񏟀5��9�+����*�/G����AƓ�\|��¨�]�����0W��v �eʙ�\����"���hCRm����0��l����X��������뾖�_��͚7��T�!�(g�4�Ug�J T���e��U(|������'�~��;'�5�;V���>����7��_]䯮̭����=�N����(��a?$F4�Tɬ���դbY�5�8#4ǔ���r�>�z���zd�1���ݷ�0f]}����>�F��NA�畒�����5W����!�v�F�w�~�PPqP���I�d��0x���A؄W�Z�䰔ù���9���Y�͉�ĩ���9���>�R���H9Y�V�u`�XUB�Z��r&��N���Ѣ[��[��x��4 Kl��g�y���}4B`�I�Z�#FZI":|<��S[F�?��Ç�ӭk_Y#ƫ����Oom��
�G������g75�̩�)���t��Q;-InV@�^X�s*5���#+pX�Y���E@$�i��&��]�7�^�O=-O���;�������l	��Wv1�_c^a����/�t�]��hU��X�x�aY�>N��0��l�w#o��^���-K�ؽ�q��W�n9�;������x/>*�0Y�A������7Au�d�Q��q,x���E�S9���ӄ��I#G�#� `��'��xr�k�N�g,����y���f|����D�[v̿�w~�V�X�������D,f��uX�ŏ�8��SO�~�G��w�����/�8��/��k��bAq����R7H"�	*5F��EBHX%��d��	���ʝG2�ظ\o��b��#�gW�`�07�Ə>$�'�� �5#���͞���&��`.�����������$��,�2p$���p�ŭ���[;��w1h�b'K]2 �\��A�gl��m2ڶ-f�	��%�����W��Hߜ�����5�"��� (���il�����~������E̝F��4(݊֠:�j���G��ލ�AǠ�mBmhԷ���hY���{:y��0fԎ@�bc-z�Dp�-\Q��0��޷��݂o��7�@C}<|w�?����bfe.�����k��Z>��ǿ%L���U�j��'�(�F���4#4�4_i˴k���^�%��u{uG�j�x}�����q��iq{z�xC��cc�q������)KAd<����aB��fH���f�6�M�-}��ԇ!FF�ae�
�2�n�R���{�2���,@�1��B+P�RV#ļ��p�Rւ����u(�9����9��J9�Z�l@Il���@� �W��@ +3��y�2��s�J��w�J�G�ܝJY��n��B�����e���%�R�Z�K�[��C�������f�Y)ǡ��EJـ�k�TҴ�)Ҵ"X/�"�.Ժ��iAcD̨*���7�B����P[k�-i
��h'^�Z�8�(D��I-u9�M�wũ�������́�	�`K}�M��{��M��0)����x�u^�jSX���@}pQ��Wb�a b[pAS8l�Ʀ�*�2G�D�-1�R/��8����.H�m� ��4��5����j�>��AQ	.	�S�H0j)�a-�lbhq��%�%.ml�k��b}0ܴ���/��7 �ii	-�I����`C[0��Բ@Z�b8��ԠL!F��E�H[S]��y9�mQ+�|Z�i$�5�ӂK���R 5 �bӢֶ�Jhv��-l�����M�M��1��� ���0��[-٥��B�A v����^�b��C�K�a�vK0X&,���6� X�9��RC�Ȭ�4f���!���!1P_{�Bu�f֑^�um!�kmD`�E��H�uLn�ҥKs
�=90s�/�E�����Y5����-�L&���T.No||@����%��g~N�����	焛�sBmr���Q	j��&�	N�#� �P�C!Ԋ���'o5B��2�u(<PʇKD7�[!�o��"��6E�:o��0����@i�BE��I0�f(�q���"�J�!:n��f�mCP�����Q6\�<�/��D{�}�@Q|s�I���_��	f)��C�\D)����1�"��|CO����d�*x���UAG"t��֬�Yq:�� ��({߬�sY���r���B���RPO���-+�;�?/���%tͩ���ô��ae_1���)Z����!k7�r�bZOg ֢��2'��Z�26��rn�B�e5�r���-��� ݵH�%�4\G�HQP���z#��:ho��rE�F�U�+���jgc��ɨ����=�rz 61	jP$��J�m�{��h6��O�RIJ���aD3]7FW#�� �rP�z�RߋZ��K�v+mɦA_�����l��?;c��RJ8�L�����R[O�B}H�����b;n�6�W}\j��C��Ζ��n��D�UC��z������]L�Ӭ�\G�� �7��k��)�в�jJ#��V4��\��|s�4�ן:E{r�s����Z)�������E@c�bZ��oq?M��D%X�rj9Z��)ȉ��@t�z���_���46A=B�	S,s�@�tX�<Kӏ�S�3�	i��˩�
�T�7�YȆ\�
�.xNG^�n�p9<I�84���Xx<o�:y���]hB�Lp1�ʁ/*�`j��ኵ�ø<h5��kͅVx"�pA�w��48�FU]8��8��z��Z'�q	L@��0�D����J���U�W���Ɨ���o��k_�k���^dC��\b�_�{.aץ�K�K,:/�g��|=��}�����q�/>Oq?ǃ>���2~��O}�_��\�Ͼs��YV:��;�Kp�64[`]���V����O�}\�&X�("��w��eGp1�*al�*��_��U�����3~�ߵ{]5��^[�{�U�JE�����;q�m=�~�1uer�=x��Q��3i.�+��������'�
&wY��L��x��p���a�������.=�v�8)s��=�5�D�'��F�܃E�=�D�aN<��3L������g&�a#*����	..va��bW��]���\�����vH;���d�E��`�=�m�k�.EcA�nT�>\*eԻp����n;������I�N��>����ݿ��K������^��6����q�ي�b��ܭLh몭�b�"na�Ϣ[�}�����M5�B�ؼ�ظѵ1w#+m4Y}�㐄�p�������C��)H&�oÚ4���c]�֎s��k���=��wc�]�]yw�yw�Uk��F����?!���pBU�7�J�e��l-���u��,Vr��hArY�}��)s���wͅ�xZ,U<f��$]��s����#8'*tI]����ua��
άp�.���H3
G����w*�r\���+sUta�4O~L�����>|�w�Ǵ�p<�W9
�Ufl�2��4���w��E��*#g4��C�-�3����.�#��80�����Y���S�T=3�D5s�x]4��ܥs�º(��3������7mBŃ�D*�����S��P�H�
�A�T�Gř�V�a�����Vh\(���Ig�#���#��\L��p�@�.,Ӈ�� Hf���"��hAtXn�K�L��3�-aZ����-}���Q�]�~�_�`��
endstream
endobj
xref
0 12
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000386 00000 n
0000000115 00000 n
0000000543 00000 n
0000000598 00000 n
0000001567 00000 n
0000001598 00000 n
0000002007 00000 n
0000002206 00000 n
0000002766 00000 n
trailer
<<
/Size 12
/Root 1 0 R
/Info 4 0 R
/ID [<EC8D9FDDD9AA39B7B9E03EBC0850DEFA> <EC8D9FDDD9AA39B7B9E03EBC0850DEFA>]
>>
startxref
13601
%%EOF
