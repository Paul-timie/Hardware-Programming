%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/ViewerPreferences <<
/DisplayDocTitle true
>>
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Title <FEFF003500300032002000420061006400200047006100740065007700610079>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20220929002114Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R]
/Count 1
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 6 0 R
>>
endobj
5 0 obj
<<
/Font 7 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Length 14
/Filter /FlateDecode
>>
stream
x�3�3T(� (1
endstream
endobj
7 0 obj
<<
>>
endobj
xref
0 8
0000000000 65535 f
0000000015 00000 n
0000000369 00000 n
0000000467 00000 n
0000000162 00000 n
0000000624 00000 n
0000000679 00000 n
0000000766 00000 n
trailer
<<
/Size 8
/Root 1 0 R
/Info 4 0 R
/ID [<803E8D51FFCECC947A7CB719A2AE7D16> <803E8D51FFCECC947A7CB719A2AE7D16>]
>>
startxref
787
%%EOF
