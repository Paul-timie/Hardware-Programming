%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20220919020034Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R 6 0 R]
/Count 2
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 7 0 R
>>
endobj
5 0 obj
<<
/Font 8 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 9 0 R
>>
endobj
7 0 obj
<<
/Length 1037
/Filter /FlateDecode
>>
stream
x��Xˮ�6��+��B�)�@Q���} ��4������);�EQv�a]�&���y�����׎:�Ib70�)pR������ݗ�����t9���]��O��c�n掩�|����]�9L����I���b���#O���H�C������i�s�I�.no���#f�&<�yy�,����g���!�F:r�O{>�	�n8�&6��dbF���8�;��g)�܉3��lKD�w�XY�-�W�&q�C�� �T�;e�f'�"`��J]M`��.��8��t��]�'T\�U�%�ќ���(>!��w���^3D�5�GR7���'�Ö(�	�Xl#����nTs�Pw�D��R:6��Y5e%�r����KH�����S��^�~;�joQ����O2/6�����o>Z&�M�+G1��2N�����&��I��L�o�,���EU�%�1�z$���]��t��s� F��HS@�;`�Ӑ��sVZJ4���[b	Va+��ΦrN7:�	�:>�����W0@�)�׉��h,�%s|6�ր�<J�9`��j�5f]��G��N%<KȞ�:9����]�-�X�++v��)�{�r:��� HSV	�ep���a�)�|���ʶ��P��G��Qf`����k��F�^���A��@��p�,�l�d��Ҽ�Ӹ8�\�v����O>�� ,m�Q��!iդJ�m�#�E"LHJ�Mϧ'��S�r8��L�S��>�KK}��0��ѭ��|?���c�Rk�WjwU	�끴ܻ؄x˅C�O@����	�(]�����WA5��Vc���S}�æ�K�suG$����[;�5�.e,��,q����e��F�C�Ĉ�مVb[N�x���|4hn��[âs.�[f��+Z��o�	|����:'5a��v�Μ�b-��&��[N���m���B^�7���p���_^��s��4����S���J���|�� 9�]�\�$�kB9�g�����튴���i��Ҵ�u��� 1#S�
endstream
endobj
8 0 obj
<<
/F1 10 0 R
>>
endobj
9 0 obj
<<
/Length 386
/Filter /FlateDecode
>>
stream
x����j�0E��
��P穑������>��B���W�]$�h���X�X��s-A��5|�rH��+���ex�	�_���6<N����Q�%L��v�!L�w@�l��@`���7���0N��_qԘ���� ����ַ�-� ַ]O*�%���-X���D�5�l_I�\ǫ#Ib���H8՟��H��x�"�D��Z$@^Z˵@�%#Q+�پH4��K��1}} *yF �t�$�*�w��ZZ�����!R�z���pD̺8�F"I�刨,�^�#�8�#B���,�e9�Ŗ��G�tG8qG�*-��^�a*�q�1��Å����Һ����X�T�	eq�c˫���&�'U3k���/��
�����
endstream
endobj
10 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 64
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600]
/FontDescriptor 11 0 R
/ToUnicode 12 0 R
>>
endobj
11 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 13 0 R
>>
endobj
12 0 obj
<<
/Length 498
/Filter /FlateDecode
>>
stream
x�]�ˎ�@E���^N#�������$y(L>���l˘��u;����.�*(��aw�%�6��1,���n�}n�9�K?d֙�o�t����<�=>nK���Ze��x�����S���_�.��p1O?��x}�Oӯp�b�l�6]8�:���Ks��z>t�v�<�������kK�v��mj�07�%d��X��~�����w��<r:�?�9Fm��ۭ#;re/`�\��%Y�r����[�����+x�,���-�5xG��;Y3{�q�mA�`�{e�|,�u,��-�����-�E��_*0���^�&��ҿ�:����&uK����_m��/���_�.�>.��L�Z3�/ѯK��l]�?|�K88��z���֧���K��I�����<���N�x��ߣ/I��K����J�?|$�c&B�Z3�/ѯ�ߏ2��2���$}.�ߋ�_З�_���#Â�M��`����i���O^�����4N8����V
endstream
endobj
13 0 obj
<<
/Length 10929
/Filter /FlateDecode
/Length1 16476
>>
stream
x��zixU����޻�����	IHR��$@ � $M�!a �D	��aUQFa��2E��8������.0n�����B*ﹷ+!a������W����9��s+�� ңV�"�f���w[\��%a����@�B�uM?q���q�R��`Ѳ�S�ߍ��!׊������2�	0F�Cö�}�������;��x����~ߢ`��c�	=�w��b��M!.�"�=�b�q�?�e8��nYS0��Re�F�bSs��Җ瑱��ˡÏ\ �ΰ/���Nc0�����OHL��]݃RR�������3,�3<o��[F��u��q�����O���|��j��wq��-E���u_變��Y���T����Ыhډނ��J�Ztzu�~�Bϣ��چ6����Q����������AAt'�x�x��y�����*��˸v�u��Ǉ��X����c@�c�c�������h�<��si`�A3�P#�[��V3���:���v�9hXXP��T�V*;	�AwA��o��z;�u_�D���t���+݇���u�j^@�iۺ���^��9ƨ�G�o2�jQ-^�v�=r��m�E�m����;Z�1�������ߢFT��#/���B�id����s8���);���6��}E���a��s�������2T%��ꑍ�ո?�+a��^�|C�msf�*+f�O�V6u��ҒI�o�N(/�;��ѣn9"oXNv�����ԔA�.g��l2btZ�Z%��`�)FpuQ�M�^����/�)���,r{�#�_���Ku�&�?"V��Tx��4WG$Yw�H):R��M�4��p��3�n�ϞV	��n��H˓i�K����\0�RE��"�%�mE�@#n�i'�'�C3Q�VE�"��v�>��^4��A��VZ䯍�M�,*Lt�|C3'F�Bڅ&P�aBDEA��t�Nl��l[�aB�3���Z���s�آ��5sFd��02x��q��@$�]X� PK���)��G��[l��r�/�o�+-B��;D�fBO�t�+��nk�Eo[u����u�[4�������"`7*��/�K�x��"��z<ڧ,�;�$b�6�2¤x�z?��_��uK���;��?u#`08�r6���|�DZ�UF�"��xI��SMz:{z������wz�d[R^��R&ֺ���������]�`ܦ���D���bGe��X��X� F�T`��;�Li3ъ����b" H5[�Qn C������%�q @FgDaFeD*���W$VԞ�3�� ��B*�H��)bs�J��U�P^I�(�"�	T]�̊dQ��ڪ�$X�i�G���\�p1�E8r_!� Z�Z�VY[qV'ւ�Չ�����	�ܕQ;���s�T9|TWfT���K�ͮ�E!$�A�q)E7�qW&F��F�)j��Id}0��
�1���R�p��ᴕ(n��'���@Fd�X(TƑz?�<Q�	�=�R8�]>W���@�� �j���.pSС��PL�/�ҋ����#RY%Ya���sEV3���0؄\��S!̌x3�27r��V�o���-���%�m�[���DTX�ŜH}1h7�^�&M��]��1׏&@�k���c�h�'w'.'�,���(�	���ݍ�Nk����ٕGM�Qy��̄�_� �<*¦A[�JIE$i:T�t|�Q	�V���Z������{�0��`�m�(�T�HB�p��g4m�h[+m�W;",�����4���a�1i:-/C����E=����0k:m����)1:�FHQ
�V�@]1��E=�i�	�
��Wm�H�%���W�V�#Ɔ ���br�B}D�Dt�ҞO���iW��b�� ��&0��&)&�Jl3]$��Si3}5�[	��*�d*�,��b���$�>�}�l��F�=fϰ��ef]f�J�Y%�T�R��Y,�H������{�&�/���������Ȱ���)L~o�N���}�[��F���&��R�!�>6Lƨqj��`���	9�$�H(v
�pE�� h4l�OcE�f�ˮ�7��|Ov��\����M�MO��KDf�K����{ �G?	���Q�������W�I�͂�a�ʗ��>4^^��r�]nǽ2Y�j�}"7�P,J�lA��1��4&�^�c@�����Alb ���aa���
v�H�&^���u���W||��͛wld��Y<p,���!����|�'�����4T$t���R:��F�Z��I��\�/�a���F�2�����|��C8�K�,�9�r\�(-f�yx�'���=���苶F����Խ£3�~J�,+��XR�g�����O�չ��)���!+s��V�.�����lҾgO��ы�,��+���-Ҁd3P�4hP�=��g���D�U��`��p���C2�k`�ۡ��D�������+x�ps<����7O���ޭ<���˙�]ow���}<�o穉k�N��k�ћo�� ��l��lT+�j�O����D1�����O�Y,�$c|0�l����x^���'%9�|I&���ǣi>�W��"@�Z�('0=��(���Ջ�ܑv�=05�m �L�3��̣�Q�Y\D6GJ�8<�,����*��v� �o_��N�慅�%��cYx�[��t�O���Ǘ�(�UM���e�?���ܭ��fT��W�嬲i��OL>��L�^Kl�EЩxXsʖb�`P��m���d�D)?�&%�Y{��X��6lmChŎ��}��3l�?�c�����DG��QSϼr�+p�^<H3�QR�Ec`Z�Y�՚��FÛ�Fė�PbԠ@e�oP`!/�����1�`G�Hx04)75k��<������[|'�Y�5Uø�{�%7��ko�?Nd����c����4�*�<�k5�m���6�b�Y+~���p�+�ϟ��G��<�_D����!סY�^�A�V�B�>�WW��|6���W�+���Y^�dy�)W�LWS�C�^?�FE���Qܲݥܻح]����Z�E���OȞ�4�E��J.�+A.��iRǲ�恱�����h����bm&Cf�Ok�#U�O�r8���s����>z���񬠻#���yT��>\��#=�6���'43��N�0�q�̰�|����xn(��>t=v��=����re۪��i�֓b��D�k�'oҏ�w��/�b�}��g�,�:��x��V�b�ɩ��a��x�`�i�}:��e���cA�Y��c���f���y��<WZ������>?+���}뭍7��?���|��Ɔ�T)3�Ao��b�Ĥ8T拋ӚL��LZ��wV�,0�-��s���m_�R�Ro62�G-f;��bp�S�lKx2����ϟ�FNy`;�'�����+�é؂u�).���|}�8bz�h�d3�������tF�r�������!��ɍ��M�O��Rb���j>�����:�1�7���j�;5mMMyfz���w_a�g �R"� c��f=�|���cb��F��G����`��X�jN8��y���F߉#rY�����>�k�#N�����Z:����0;�2�E�������N�����T�&��|����j4�!R`M�������F<O�:?��lׇ�0����/���/a�?�}��� � ��
���)+!^o�F	I�q��cb�$c�3�����j4ƐO�b�!��'����v-4��&\����,R@g��?~���K��ǋG6�z��Gv��"W�g��_���<�ų��g�@�v#�c��Glx���_��|��Q�t�JX������ŐOo4:�;�����FA���ݞ��U�&�kR�������=��2�o�
���7�jI=o���g;��|�����>c���'0�'ï~u��o�\����ZK�LaN���k�mK����g/F�g>���=u�u��Eu������$I;,���xp��}��F3�w���6��ObT���,�1��%F/`-ֳc4���V�����6Oŧ�m����'�D��y��FE�>�"�`V�b�������V��G����D�6�&s@r�J�4��OFf��l1�|Fp��ºp���.�I�YŐ��+�;n!$QP��0��"BbX� �+wD��,���zb�h\hT�d̕\��O�(��Aظvۜ����37M��ޥ����u���O>��n~���c��YV�`��Q��-\�<h8p��F�8�!X�f��Xsx�	�EI*��6 9&�lֆ|fN@	}yܳ��(|�G���r�7{�Ў�m��b:l�N~t��[���b�ز�Ӎ+��
�y��}���s���S߱dQ���)ל�,�u�Xà�Se��f�1Z�f6�T�����`ɮ���e9���}9��5`䁴�g�vY�+qm�^���
�/ߟ�����
u�����N���{Vn��?������
�/���?�ͩ����������>�U��Jih|��j��ԪI������fKL4�|����6-p�}���z�o�"����%B��(���En+xo��\ɒ/����.l��캉��G�YW��Z^8}[�Ah�����<��ɬ��=$Ϛ}��.�4Э���\�cX�9��(9�*��*Hg����Z �N��\0ǹs!h��1�Ε�<)u�.�ź�G��J����̃o`���w]��E[��=�j��W��i�>|5�V]��q�Xr8�S�������&�s:�����)��b�Z�0��$J���=�F@���fSӬ��z���| ��e%����L�v^<j�N�<��vMA�;�$�۬��?^�{Qlޡ���?~z%J�s �A���)����^��U��ҝz� �uBS�c&V[F���G�7twԿ(4k!���N�������f֠�N��p����;v�޽��6�~x*�A�.ݝK�+�}�ӛ��'�Z�9�yij��I��G����x��1�g���K^ǠB)U�q<����»�/Ǹc,���q�ׁ ނ����G�ܗ��,҃!� �v�`��c����~}_tm���l5�"�ں���a�p@V8Z+@�Q0�Y���|:��M F�=�k4��+Cd��r.�A�-�L�FzQ[a�۵���x��1�K�~N����^���5w��Pqp3b�����kֽ#����?���?����(��	�K|O���4	�f��^�#ƮFƟ��9J�Bӓ�������z찒ȍ{z١g��]ӷ/��dB�Ds������&�9�N�3!D\��Q
oOIMKM#1���M�M�c'�xy���|�����x���ټ�pc6^suX5U7�����u����p��ay�a�C>f�t�<�����IuuT_ڨm���H	����OК!�!y0��1�x.�Ġ@���v��< ��L�K�OXx�/��I>�]�p>��>���3�c������ڍ4$:�Ju֎�Q���K4�e�0�)�	ք*��
���F���"R%3�ݬ��`�DE�K���p��V��͛k�/]���v|e��ȗ�n=��9�P�:�|�x�-pG��_�j�\-�j�S����(9 ��P��1V�M�����֮2��8�	!�<���Oi�[�T��q����a��<�0=�O��om;#�ە�s0 8� ��_-.%����e��^�a�.��	����{@���c'&� �>��������4l;*+�u�,aN��U4/�Lzd�\��6�2���X�S�ȡoz��\�.�":�˩���� ���~������%�v��ˏ>϶��Fc��}tR��0��"�b��&��)�l�z��b.�Y��P惐ZI�r��?7!����͋Z������ޝ�{�cw���L�[o%��A�y�������f���[��_���c��V�%&5Y1�����&k���*hX�o����Vk\�	Y�����MXJ����nsoD�U7�V+5=[�rB9-�+h5f���BR��uɓ�<�E��c����n�$cxp�aN�vf�b}�o|X��K�R�Tɢc��4��XԹ�7e;��r7��{m�w�v�x�� K�r�xVQ8F��k�W�,7�U�\E��#F���zSV�3/=�;�]_>�GW�(������<��z=k�XX��p�=c��e�-����岅�Cd�x�L=B4f�w��{[n�Ɓ���Q/f��~�}U~��	��߯�����=�
���8���_��K��N�z�=sV�J���� �+iY�*{��<��x�+��xō��iP�����0�Ց3,#���0k�bV�b�>�c^�BU>��5/XW�#"5���b�x�����]�^��d�|�vz��\ vdG.��%��1h��_�3�L1Hkg�e��_:OMLs��ѽ������x��lFż ��qs��k^���G�޷u�2f����uGN�~�^���[]�ϝ�����~?��oo0�3��$tUN_���pj�X`auHWQCߴ�WuR�ȑ���H�<��)<F~�p���۹z΁��GY�rv�#%0��8^�����Q���`7 �\'�6���韗�ߋ5��)��ǺҵL~�C.��&I�?�1 I�P���f�ǳ�b�o��x��T�$�L`����x��CɹE��\�I�b�Đ�ݖ��&s\�����IG�"��xf����zp��o���\汸�w�_��YV�nyUan�xץ�jY�쭼�mRP�8��+["���GcJ��w���d=A6� 9%�9O,�7�\�3V��_<�섨p�vн:�E=߱�3%=�q�jU>�Z�|d�?s�^�$y��5��M�k�:�_?�!��/�>%�-����Ooa���-����@����{�y�������S<���D��ڵ���DuG�)>�\[勋c��*�N���0kON�cy�_:J�!J�+��
$b1�8Qn�W�	hPc�z�콽O�������!<	��3�÷����׮φ��l'�k�r���Jiz>F �Ͱ��#��$��Q��g�zN��:A�u�����}�]�z�yu��5���}��������Ͳ_���k8=���ڍ섮¯��/��(E2k#H�b5�XVC\��=Md��=�17���W?>���S�����}{cv���w����vXg��gKYY�V�u`�*.^��W%&��N��Ѣk�ݯct<l<4��m��!ozL�'���'�v��4�z����V� �@�����Qi{�p��\W�u�k��X5�4������1�S��v��{�Y��gW͌g��.��R?%I.V@��|vB5ϩԜ:F�4��a5gт�����~�a���!i���y�:<��<rFn�ם��ȓϰ��Zѕό�z�y������t��^��hU��X�x�aY�>F��0*�F�Cyb�^-��/�������'�9�{�����Cx7>&2��A��������fB<v�#�sHF�NǱ�AU�q���`�O&K�;����@Ba��y��ݯ���X�r��H���ȕ��m�����i�,� "�ٟ���Nd1��4��¶<���ƞ=ot������o��O�*��z��?�ȥ>+?����(�X�Đ����pd���灈�g�{�IԱ3(�+�Y��o̔n尊�`��g��&nw��XN�8�!�:���e�7a��8��ÐIя����n�}�Zɧ�����_��[��h˖��'�Y�>0�Q��C���Z��5��q>
���ߜ-�b����0jl�������@�g_����!�h|B�w�?�[%�>F���BPX)��-�FX7,�D���7a�x�+x����z�zB~X~�q*����̟��r,���Z�/J̄�^�����+��~���2���qF����	˟����k�,�}������y�ޮ���K'��_<1w��S�tZ�jЋ����v�M�}��Cyڀ���݌���U�9hoCG����wAX��S
�{�8	����h*�u�a�&9��3A+X�6��� m������pL���0W�:v'���5s�y-���
�������o�3�[�����4j"Z��X�B����l]��^�����迎q���=�3�p��#g,4�62~nbL�f�n�qʙ�(��� �F�CZ~�5��Ho2n����^^bd�Vf�P@)��7-R��y@)�ȀU���V�*��+e5���F�d �����gNV�:��t��'|�R�Ay�V)P�O��4P����2Fɠt�2��[)�h87L)s0&��y��ݫ�(�P�*t�{E)�Q:P)kP�g��e��U�:t�����ݮ1+��P�X)�p͟4��j�Z�/���57,���5��ܜa9�m���EqB��)��7��n�+N��p�8��&��a~ :V�lN,hY�o�	4��š�Mn��4�H97+''�s��!�/��������_����D�́�p�Ŋ��,��4�Ec�8�w�Ժ��� m�	4��08�:�47�jj�PV/�}XQ,	����p l,�� P6!�jhd�K�j�ť��X5,h�������D���j�K ����k���!cH��b��&k_77��-Zb[�S烜�6��	���tJ`龬j�Au�X�aqSsp	%th��9h|�Z���Ea�U�o�� ۀw5!�����oZ��l
 ��n+�1ȋ�4\�$����I-,uLċ��_�%�����p��>t��05(�kka���`M�b",�u��8Ms���� eq(�>n���t��,�"�O@����𲦀"�fe�RЁF"�*d�����&�����b�z��� 664�CY��EY���S���5�n �� '�j���~(���ل���'��UD��:޹���-��`T��|M�r3�"O?�D�(��	�Gh�P��PQLggBi"̯�0o>���+������v�z��u�`N zj����!�r�L��m��r���<?;�6 $��8L{��)忂� l���	���B���Z
�����tT�I����?�q*`���5T�=#k(l�Q�A(�+�\�n���y=k����kE9�n	�9���z��@=��+�3��J��	?�5w=-�)Ok)�a�����s�/���~E6�TrKJ�(����3D�6�~�j�RK8Rw"嚟� *����ck�}��)ֶx�:_����:�{�OfEy:�K]����&�Au���n3]���R"�	P*I�O�>�XD�F骧z�R(RS�{�V����n�-C!�k�8�(\�a��ҟ��^_-%�YD����H���m�^N�Q�L�/�>�W�R����f-�6�?��&�`R�j��{TÂ0��J1jYQ������Ae^�Ma����R�6��^fu�E�����(֓�М�=���D9��J�{iY4�*~����Z�Xr�$���R�Ѥ�W�xb;7{�a�o�M��jc�Ô��e]��
J��4�d7����Ƨ�rȫ&�
<]y��3�9q���<��T�Rx���h,�10~4�o�:y���Z�h|�Lp3�΂*ƹ�j[�Ꮆ�y9�j�'�;ښ��F"<����"-ip�!�*:��Cc�+�E��loƅ ��� � P ����q҂
ԅ�+Kw~�Mw��;�yś��tiǥ�����M�������y��r�2�.H�yo��_�:��r��/���/�/>�:��c�s����s^�s�;{���yFx�y�ǰ���k��cي�c?��l�'h�;�"r�ay�aYvT7��R��R9���R!~R�I�'�O8�'�=��Y�z�����'N���R�MǱx<�x�q��x�q�x�y��>�,x�౳���R�bGNGYGSGkO�0%uX{MG�x��H����p�0c|1���/�8F��W�l�l�0�Hg��}0� ��@� �y�L����̎�q���1�c��b����7�0Iv\��z{�v���R����:s�J[����I^B��1���Ԗ1Ν�5���My{q��^�|4��i�rpˉ-��e�0��ő��k|$���GV>r���2֣ �K"���T�C��γ�q�f�ܜ��	n^��A�L��M,�Ķ).�+n���L�P�!���Y����׳�z��k:�u�
ʁ���ĺC���()He&�w��T烓�8׮�\s�����;�Ǧ���r�cs��+Wci�F��|��\�p'ชxO\���V �j諂�h�9�:�L�҂�&y��.v�������Z*x�Vp�,h��p����Gq<�;��:�����Z) N/Kt^��=�����╦��{�-�gKq�w���[�,����|<	�1+��6�z�Y�e/��ű�^�ȵW���k�`��0�WRb��i�7VWB�o�6N5���g��FU>�]6�AN�t`w���3�32J:T��K"��9�6�RN�Ҵ�amU̞Sَ�F��6��%����H� _I�
)�B�4�݁
|�p(ܒ��R���p޴B{�F=&�
�CJ̀Z8��>3B���d,��!�0)�°�f�0���GJ�4/���huL�(-���E)�`�WB����n
endstream
endobj
xref
0 14
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000392 00000 n
0000000115 00000 n
0000000549 00000 n
0000000604 00000 n
0000000761 00000 n
0000001873 00000 n
0000001905 00000 n
0000002365 00000 n
0000002788 00000 n
0000002988 00000 n
0000003561 00000 n
trailer
<<
/Size 14
/Root 1 0 R
/Info 4 0 R
/ID [<BE54147345785CD1949AA1D0528DC8C8> <BE54147345785CD1949AA1D0528DC8C8>]
>>
startxref
14582
%%EOF
