%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20220929002116Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R 6 0 R]
/Count 2
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 7 0 R
>>
endobj
5 0 obj
<<
/Font 8 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 9 0 R
>>
endobj
7 0 obj
<<
/Length 1121
/Filter /FlateDecode
>>
stream
x��Xˮ�6��+���Iɲ������� ������!�ܹ�)�` \_[����e�S����u�w<vQ�"u1m���u�����Ʒ��!��E�ԝ��~]�#ם�����?~?�{X·/E�(�C�$v�npэ.��qU��=����f\��%hH\tq}�H}�c�
���L��1	y
4ؕ�l6��FJv����XU]�p([H?�t�~�ꪸ0�Zwt�Zy��8hZ�Y�݌WO��w��/DvU�>�]��=#|���-��V89y�{��&�����ʾ��@	�|�43�{7> ����\+D�j���ͮ-
�����C�zF���S��lTu�Pv�i��ťn�
��hJ&�Ƴܖ�����u��RU�C/E�M��E�aW55vJ�O���%���d����I~oM�+g��je��$�!U��1�%i�.?�����,,"�"D����L湡&�2��`��*�&���%*w�./�mU �[+� 9aV��Kb�tE���q��
�˝]R��'/*�
��L�]�{��}s�Lg�x3�eӱy�rr�UhB%f�CD��w�-<[��Ker����*:��:�o��`I��f�X�1�d��Y�N�2l[�lL��(��o���U��P��[���W`�F�I%�_��Z�����ykی,y�DR�*
�!��\����\�L���z�CA�k���#�=خ2]�_��|�DX��H���&����?�I\��S��qul��G����1����vX�̟��=�3��;���ZN�Ygk���l��!5	
���*#ΫQg�W+�*��(���t[��U�A�HaF�'�Ӻ)k�k6��B~�+M�:p�$c�V�}6$ΏZ-H�}���hh�z<�@U8.?�<�0C�%y.h�U0c~ȼ,�ZF�%�!Ew/d/��}���I��-��׏E�p?�_@rDc��.C!;�����B?�s�5z�~@*�E��Ok����K�$��S������£�x��۟����C֬�99�7� �� �G���@�Հ���V�2�w ��D�ujG�x��r�Q=�����C�4�|3d_ >8K�|�� �
endstream
endobj
8 0 obj
<<
/F1 10 0 R
>>
endobj
9 0 obj
<<
/Length 327
/Filter /FlateDecode
>>
stream
x��T�j�@��+���v�}C)$��0���ͥ�_9��`{ݲ	�^iF324���MAA���D:R!����<ܨ���������:��^'�?�ێA��w��[��&[�	�p���R0������}��CN�Z`���Ъ氚+N�R'���3��k� ����YlI��F�䰑����<��8I�r��C�
� Ol��z���:8��|YPU���*.��:[QcÜ8���(77^~.�ڊ�j+�Ή#ƌU���!��E�Z� �*ђY�`\�2k�yHU�X4+�5fu~Ϊ��w&O�/�6�\��&�Jgg��R��}�(�W춮'
endstream
endobj
10 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 65
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600]
/FontDescriptor 11 0 R
/ToUnicode 12 0 R
>>
endobj
11 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 13 0 R
>>
endobj
12 0 obj
<<
/Length 502
/Filter /FlateDecode
>>
stream
x�]�ˎ�@E�|��b����d!y�X�"œ��v�b@/���[��HY�:�T�N�)g�aw�5��L�ѯ�y��ߦ�����/Ø��C�Ɠ~w�vN��{|�V=��i�I����m]�Ӷ�N�S�}]z��%}����x��_���5͓�N{u>����3�z>���>�Cʿ����S�gC�n��mn;����'�<���~_'~��{VL9����BM�s��[re'`�\��Y�K�J�+����ʘW�VY��7�/��+�����d�ٳ�lr���)�_�c�/�c�o�o�/Z��������_л������iL���+���C�&��[�G/��e��\K�n6�#����}�?�m�	���m�?�l�_j}�Z����ҿ������wC�y
���1[��C_����������п�L$�?zO�J��_�_��L�L�n�u���7�[�t�=���7�,q+�6��?�v�e	��˯;��F���a�fd��7�l�
endstream
endobj
13 0 obj
<<
/Length 11054
/Filter /FlateDecode
/Length1 16648
>>
stream
x��zy|SU��9w���IW�B[�+A����BY
�ЀІ6����&� #���*�(� n� )�K����8���3����63����Bo��ܖ�q�~��������{��<�ٟ����� I��M^��u!l�^k9�/ ļT�4�Gﾎ�!�+��ֲw�݋����b]�_��e� �auа�s� ��PP�0|��1O���nV���Y�e��B�}M��&��C]l�/��,
�k�6C��(UF�����h����*�o@�_m>��CQ u��xA��hu���d�XmvGl\|BbR�d�������6p���̬�!���yÆ�1b䝣F�ɗƢ��/�,��/BvTE�}.n$��%u]"��K]�Ѳ<S���u��
z�G���PzX�Z�@ϡ�>�O�3�E��@;�F4�߂=p���VT��W�{Q݇��ux��\܊YT��h%j��K�6�y"���7�ݏәm��6�1�_�G��Q��ϣ��A�oУ���<��u��*f"4�kOF���h.hX=`��T�V*;�A�CiQ�~��6���C��zt/���)݇���u�n^BGh����>��9��;�@��g|jP^�v��r����E�m����;Z�1����
��ߢF4�C^��OM���x3���2p��� \S.v62u�i���\%��#�����o���RX��!�;*q�W�?�x膤�f��U�O/�6�t��IK&�/��[T8�`��?f��;G��c���!9�Y��RS����q6��h��i5j��s,�Q��UE6E4{��"��83C,��+��(r{�"�_���Ku�&�?"V��Tx�{5WE$Y{�H):R��M�(4�,�#�
�b;�5���>1r��'�2�J+1Pq�`Ŋ`+E���Z�� Gܦӎs�h33P�VE�"�Mmx�L����mRǐea�E��H�Ԋ��D�˗�1>bp�.4����"*
R�'���b[FG�v�W���q��ﮈ�~���������#�܅�A˾���"�¢H:�Z2�g��[K��br���!؎��-~�EH1}�H1��i.r%z�֭�^��m�j��w��s�&wk�^��T�F� �������_�TU�G���{��D�SgWD��X���]w$��=cJ�]7� q��.!��v	̓J�ejE�.�y������0U�����^NzZ�{z�W���%e�.e|��(��i�ҵ�0�m��Ot�[-fqD�����5�b�O"���@nȔV����.'��f�8�`�"wQ��]\ D tqzT�WD�B(H~�cEm9�0�_�/�̌d��"6wAw	ZE�et�2-bAU�ʬHv�+����0���Zqy�.�_��!����q e�E�5�gUb�]�X��H>��]��
��H��GeezEI��dꬊ;D��RtwEb`D��+�D�M� z��.ψ*E�	N[���+p"�hD�E�Be���qW�M U�3�8��sE���Eea��&D-��3j��qŴ��2��X��}�:1"�V���P*+Ġ4Wx5�O���L���B̈7=�7q#w�zO�������b��]R�J���0AD��;̉��v��M��T�[�$�(s�H�=���]V1��{��ed-*�%�23�����کm^[6��	b���+3�WU�k }�Dp��!���TDR!��AEM�'�j��m���v�h�����v&�f�.�J�=\�G��A�:��B��Ն�$-/�%��gb��6L�C˫�j0zY�cpb̚F��qK�FJ��h�Rõ巖.�U��4���
��W��R$�AY�k��eC`|q�� ��c AѺ�������h�@�U �؁az�4��̮p�J�	g[M�	�|`TZM_fr+��d�@�Bɒ^@*�jO���s���<b��c���]f�ev�`��2Le�tZ����jx2~�}�i8�A�ѫ�l�1ʞ�N���y.;�����w�&��]����,�@)�l2	*U��c��d`������J��l���#H��Ra�.�A�
�F�V�4V��nF���ʹs���d�#(�!�=������6<�q��lr�VUv�g��#�gG�z\>,�(���{S~3���}�U��G���\ƴ�mc�}P&�_���&#�E%�E�#��k��>�����X�����{Q�X�Lа�CS����(q�o\��?;�v��k�رe˖]��dX�<�8��_�_��������H9��5�v*��;��@(��d�Z�I���\�/�a���F�2�����|��C(ԃ|,�8Cr\�(.f�yh�'���=���苶F�됱Ҕ}��ӿnr�L+30X��v��������Χٲ��ȩ�SU�`ց�wf���{;7B��^�gr\)P̍��%��8�AR쉥>��U'2�R� �<�z�wz/�)]����d&�m_r��}_�sG�C����z����ܾz��/c�w�Ӯ~J����a��:��(��g���Go�CR��]�폲Q�42��`Q���b���b8�g�蓌�����W��y���(�%���R���x^�'� Q�J�"�@�l��X�#OT.Rr��w��4�25ϔ2<��G�fq�)�c�h�20�EnR���ق0�m�S��[���iOd�o���?U[��\���T5�ꛖ.8���;M�0����ҩ��ON:�TO�VCt�e��x�sʖb	cP��m���d�D)?�6!�]z��X�0*6lM}h��W����3l�?�g��}�Ȏ΍DF��S�?ݙk�\���)Ѣ10�ɬ�j�v�A��MZ#�K}(1�P �ٷ0����iy���{�#v8<����5e}�E܁ճU����S�L�a��!\v��Yˍ�.�$�����1�B�a�dX�5���v���f�G���DX��/�t�#�H��.�=@�y����Li�� V�U!Vë+}N>�g����+��!�<�r�<����A����!K�A#����(f��R�=��΁����E;�YOʞ�4�E��
.�+A.��R:ǲ��c5�ٙ3$�hK)���L��R��`G�R���p���	'��y�P��mYAv�'���Gm���Æ{@4l�U�O2hf��=��n����!/����7���B&��^>tm{p�2O��|�W�h]_2�yz�̂[Kĺz�f���7���K����|���C��G�=���jP%9uz=�k��F��̧Cjؖڈ8D��+#�/7����z���<v��x����y�u���ooڴ�M��AGGt͇�VxAol(M�2��T�V�*�ML�C���8����dҲ����U�i� h�uȞ3�o{�R�Z�ᱷ(j1�1X���0G�S��$�x��7r��<S������&e.�b�a���|>p�	\L�����A�� �˵;bV+3�g5���6<z�;5�C��ɍ��M5O��Jb���|n�C�u��6�7�e�ym�խMM�yfz��Nv]c�ÚäD��f3:b�z��5���,��� f��e}��5�c��9�H�V�O�y�ȥ�����{~���&� ��3<eb�uY�2��<�C�����j����b�c*�	p�Jg�9_�a3D
�)5���\@>�܄���x\�'W����]&"�w�E�Q���Ǎo����� S �!�A"�.e%��-�(!��1�qLL�d�w�3v��Fc�4*����|�9��[f�Bé�h��Wd�2�M���o�_A]?^>�q��<�{�V��"����W��x�%?#?��c��˟�?b�S?�����Ӹ̍*�;T��Ϣ��K4 �(�|z��i�e<d�j�2
Z�hd����Ϯb5!_��EŨTd��9}��י+d&�o8��2�
z��a��;��|�����6����'2O�_�����?��{Ūm�Z&��̜���׬ߑ����Z���}�O�{��K�7*���`3����EI�<l���x0����~���;|�=�'1*�[@~F=����K 7$�l[���Y�U8���yv���o�p�P�����n���l�ʀU.��!�޵���ycL���鏮�z���\�-��'f��ս���툄������2Fm���RQ.Z ���gj�b���cb2{Țg(D�f��:Y���i�)�S�|))���$��9�"n�e�t�=;�F�$`�6��`��`?d'ɘlŞ�oqN���ɼ?������oZ|��ugZ�V��t͊�׵.ǜ{�Ƶ;�?���������K|�i��
�S�{_rp�6�]�����2�徕��ll%|�
|Y zm �d�^�Z�g�hR	!H�V �{�c���v;O0����0����)���[�j�����99�uU����P9 qa	�{0Z,�M ��/9Y%�@�:=#�b��C>#�q�ba]���\ .��j��!�k*�G=���h�~ݣ��t ����74��<��"Q����g�B���Ƶ;f���Λ�y��.yL����^|j�����ճ�O�z`i���;G�ݵ`ɲ�����/,�$q�ð秀ƙ@cʐ�˪t�""��Ԫ�O-0@�>��$�)2�M+xP.SN;��7�Nv3�jgE��b�(����l��2i��a�_�Vs�qF�
3:�ҧ��f�q��0�$"�VΙ��-M��z`��t�.֍=l�Pⴭ��ֽ�����u��m���ȫ����sG�>�}�zT�W^%�W*����*�)&�`�Ʊ	�Ng��wuHz��تV;��AA��C����o��XP�n65�
��cu��cpj�>���Ϯ{�2��}��=;!��_ؚ55���d}'���N�/�y�gm�_�t<�� � �KE���*�i���U��:���"愦F�&$8L���h�9h�#j#�%蠙��D��D�IDK�e�f'Nf���?�vY���6M��L䃄=���|Wv��g6O�yOZ��9cʋҔ���e�=��
[��΁����x0�:J�*��N����m�x��c�}P��q- �-��~N>y��g	�1�=� na����2&�n��i7��E76mY�V*2���+.|�2��R�X�2���=�j7 �X�өMl���G�Ii���E%>s��7�m�n Z4z��&;wȞ���k�>3�a^pB�_��~tÚ����R}%Ķq̰��gnX�3��qç���Wz�]��1�r������i�v;�vG�]��?��as	)�;�4��X�툒��yf��縑��v.��fB7F�9mg������t7��� ��@��Rx{JjZj��͎XGlZlZ;�˛��`���#g1���c�&��M^͍�tÕ�j*/o
G�?�V65M�
|G�$=BI���ꯏg��*_�~���$�
� �֞��od�s�,MH��dҲ�^2,B��&s\�����	ǒ"��zn삇�^7m�x!�Dܖ_�_��^Z�~Yeannצ�\���[q��<���q���[#���G�J��w��i���S t�C�^)�7b ��ݶx�wm����Ny�_:�h.������7&������
����y��_���5K����W�9u�a��˲o��ow��p��O�����|%�^^)M���Z�@Έ��90�Q��g�z�(� `b�I�=��9RlOJ���P�k����Jg3s�oO�[d=���!u���.��v;����.D�[���Q2*����[9��NQgM�&T��V��,4RO���
U~�H�H $p"d��d����$��ɵ�W���N|m����W�o?��1�p�&�z/�m0�ǖ=o9�?�g�\%�l�O��1rV<��)�c�V�Vg��6�]e,�q*"ae�`�嬵����X�}숆���=BL���;[��vfw���E���Z4TJ /)0-�h�N��\9%���m��}>B�u��NLNG��}$Oy��C�i�v�^�k_��9ݓ+U��
+YI�L�#"��ƛ���V+}jV�P�ߓ��29601."��j�l1��rɟ��z
������{��ٶ_���)�E��;/?J�^$�d��&��0)�l#��v��\� ������w�(�o�FV��+/j���-��ޔg3����*�3%o��t����-a�3��cz�{��	�NJ�A��XmȖ��d��j�VY��-���a�����ָ8$��\�����I���D�[�]z�N��jB=nUQk��A��*�\��KI���O=��o6�O�,ys�w]�I����V���7?��܂��������LTtJ�R%�
c���4�#ڃ-��>Z�3�yR.�r�n�����I`A˝�6"W�g�c�:=؉q��&nT�ris��v�-YuKμ�x�����?��]�������PL����AcaYN��:���)l��[��S��^�5�y3�Ѹ���Xh�uJ	�Fd��ǐ��v�}M~��)��߯�����|�m~���|�/z����&t�Ȟ;/n!�qгA��+VҲ�h��@0J��I �F� ���Q�h;O��1QF`�:r�g�Sp%f���A��Y,�c̫T�ҧb����j�u4D�FNB`3v��y���S���>��T��|��;�.�:<BJ@T`P5}�V����!]%D5����P�S9T$�`���7�g�(�MX�Ʒ;wr1ԗ�*�q֢���H	Dk*�8A�ṝ������Jzzz�Dv䲺����a�|&zrzc5��s��]��w=�풆�ac��c��
ė���IUUT.��'��y��#�p���Qȹ)��.�bvCT8s'�c-؀Zzfc'�D&zZ��*}��V�H��3�D��f�ˈ5�ǡg0\���~��\�?�������SO<���'���Z<O�='�g��o�K�_Q�ob��(|�!6���v-�&!Q��uM��1��V����:�ҧө9�#�`�D 5(���!>1E�"J~�"��D�Æ�M���?j���B/����i\^�h��1>��8�'��x�|䎿ޔ����`��zm\��s��R�99Y�L-�6 �yo�#���hY���h�뱙��5*�u���V.BuxN�{R��8�9c�����OV��o?�$c�5�_v ��'�9����'��P���؎O~(c�����8�_ߘ]y��-��-)��ٽ���`?D_�(E2k#l�b5�XV��}�EM��ă vG���/n^��Ԣ'�^u-��E�م7���쇬���Js˳�[z�h���'hͥ>bqy�������;U��ډ�0�~,x�+ l��)~ap���C�E�����M��Ĩ��Yus���>�R;�'fIYY�V�u`XU\�Z�JL`�*>2_�E�H������h|&��!ozd�+Ԉ�9*��F�]��b6�Jޡc(�?��<"m����J��y}�����?����k�G���{�+ϬoH�U9#���x ��Q�&I.V@�Ì����TjN�GVచ�hA��I�S������!�n��0�x�9y���*�?�?�'�cܹ�3����:�].���#�.�5�
s�t�3,��Ǩ�� tf���yb�� .QW]�~�g�S�k��.9�[����C�Y|B.d2�<?�y���{f@lt?�d�Q��q,X\���E\�r�����%֝J���{@���;Nv���';�3��\x�>)��vIG�/�����Z���|���3��X�&&�㰰����xs��7;������w]�~�`=~��䉔va�$7��*u�$r���Rc�q�/�+H{��� �2 z������8k���f?��<;���������4v�
n&{���ҝV,�����\�����q|�IG18���\��p�J�т#�}�G��@���M� x]�	���ي�[e�u+���{v�Gz���a > �\�W%>��́��.����e��즋�3kY��(�V��xmH�1'Hs;U��ip��,���O>!E���s'V~�9BcQ2�hː�f�͑�%��'#���n&Q�)]Q���{*���c����=n����!��~����0��u>��o�����b�Z�'C�^�
U��Q�c�A���0����r�5�-P�
#���+��ފ�a�s�C��G{�"�4"�= �4zWu݀x�V؎6�;X��x.����p��h|v����p+�1�Z&�\gk���\.���|���T�+lS�TcT��OԒ���F������}R��N����}������_�#Ɣ��Ŭ�yېlXmh7�d�a�f��ę��jMϛ:L��&�B��>���P6�R�c��Gz�qcg��##԰2K�J��\�A)s0f�R�=��(?��UhjS�jd���5� b-k!���u(�����~�R�Ay�V)P�O��4P;���2Fɠ�2��[)�h(7D)s0&��y��=��(�R�*t�;���h H)kP�'��e��U�:t�����ݭ1+��@�P)�P͟
��ׇ�j��/V��6�ϯ����9CrĻ���q\��)������n�+N��p�8��:kb��@t�8)�������<6Th�	4���mn��4�H97+''�s���!�/���5����{�`m_$�����P8����byVY�X�â��F��3qJmm}u�6V��~��5ׇj��j���{��,X'���@(�X��Z�ٸ�P}c C\RW_]'.�Ě@�~~#t�[*��%B�v��\@ô�@ms TW�8_�Cb(�\_���u�0���@�����аض�	��>-�ב����Ɂ%�����a���M�����Pus ���k����� �������C�,@��ߘY��9� dg�5��@@/J�P�aq DG75!�jL����{Ȗj�̀fM�.�޵��0L����;,X�h!a�:܍���9}M�0@Yʪ��Ffg/Y�$˯�ؓ���/��)����@Y�0d���oe2�D����&����b�x��,d�o
��B�Y����S�Q!��]&�N � n?��P�ׄ���'��UD�u�sQ���QA�o��"�f�E�~
7�Q8�q�Gh�P��`QLgg@i<̯a�<��WD��;H���� ��h,
�� ���"ʄ��!�r���i��r��N��f�2�z�$R�i�r!��h���%J�0.@��� ��P�v9�(��J�LB�0]�����3+N�ka~5�a��j
��Br�u
= ��)5t^��B��R�祢�b���9���z��@=��+J3c�@#�z,l��u��4����5*��̉������+�i��[�`�XY�P��>Ct�FXC����Z����ކ�H��<��}!���jho��RE�����S�i	�κ���YQ�N��W�龴�JP�"�dU����E3)��~KR�S�3�Q�ꨜ�)�
���n��(�$k7іL�5�(\��L�b�z���p������b[Cۂ=�&����;n�6�.�RɋR��B��7����	+�)F5���=*aA���r1�YQ������Ae^�Ma��TS�6��^fv�E����T+ړ����=���D)�[K�{pY8NT�@c��-��ݜ(k4�Z�&E~�
��� ݹ�z���ܶ��4�C=L�	QZf�=̇�)���h,M/���g����r�I�OS�3�tdCN\o'�� d;�x"�I�h4���(?�wB������-N46E&�zgA��\0�-��pG[���h5��m͆Vx#�UpCO��48�0F��8��h��xu9�ƚq!  � 0 ��@��C}�4�u��J:��t��;�y͛��|eוCW����W�SW���y��j�*�.I��Eo��_�:��b���/���/p��?�:��a�3����^��]8��.x�y/x�'���X�*�G���G����џ���� ��m���'�m�Q)�"g��2���g�I��I�'-�D>ጟ���g��7V���:�_/Mu6���ɜ�'٦�-'�	�	&�D����C'Ο��Lu��9��M�-�<��'��:�k:�ţ�G[�F�r-G"G���/_}�m�1R��bgKdK��D:"�G��C����#����d��`v��;������(`�&�E�Y؅I��ҝU;�v�OlKu�ڛ���.mg ���9���6�����Q��c5���Ky{q�4���xb�Ӹ���S[Yik�!^i�#z���X�c���x��c��U�GA��D�э��Gʺ����-ع%{ܲb�6�6��Y����$��)g3ec���F6g6npn���JLV��$�"�9p�]Xw8V�#��d�_��\7a�s���5�r������06=$>���� ^�
K�4zo��j�;Ǖ�{��U�\ �VA_%�Ǻ.`�ag��$�5�;wV��n��lxς�5�R�c���eA��GG9�,>��q��<���؁�v��R ��D�թ]Sij�^ij�@�{���D<���Y�-v���Di� ���}܇������i��Xl/w�����Xn�5�3�i�+)���4�+�+��јm�b7����|h�jd�����<n�[ڦ���������D4��#xm$��<���"��*�5���M��7nD�J"�e��~��H$Rh���_��B�PxQz��J1����ax�
��w_�Tpz()-0j��E��
uO$c��` k
���!~^0�,
�q�i!xt/	������΅) !ť���(���������c
endstream
endobj
xref
0 14
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000392 00000 n
0000000115 00000 n
0000000549 00000 n
0000000604 00000 n
0000000761 00000 n
0000001957 00000 n
0000001989 00000 n
0000002390 00000 n
0000002817 00000 n
0000003017 00000 n
0000003594 00000 n
trailer
<<
/Size 14
/Root 1 0 R
/Info 4 0 R
/ID [<C07FEEBEFC5F355E795E070176BF5684> <C07FEEBEFC5F355E795E070176BF5684>]
>>
startxref
14740
%%EOF
