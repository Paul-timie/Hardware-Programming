%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20221103023811Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R 6 0 R]
/Count 2
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 7 0 R
>>
endobj
5 0 obj
<<
/Font 8 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 9 0 R
>>
endobj
7 0 obj
<<
/Length 1043
/Filter /FlateDecode
>>
stream
x��WɊ9��W�هEHJI0�z7�x�����U�d�T�r7#:�sы�E����{��3���n �S�.����������֏���z�C��C���:2��˟�~�����e�^>VM"���X�7�	&�dF�M�z��L�>��k;W]������ 5����n�A�eɑ����SG��WG�'�bSt0u�!l��g��4>�n���k.Gʹ�%8��>Z��a�bZi�pX${_ೀ}hi*�Bݝ,�t� �!�y�쀢�JzmpѪpp���^]wʮ�*��ps���(8��$ۻ���^�誀�p��f�6�d��H��
C&�B��?���F57u���ݥfl��Z5��A�q���G��D?0MMa���귀�� �G-Hj��ͫ?�x�	nރ�Ub��W�$�Ip�P
�"7��I0.�{��%	�@�њi��Kxn�j`m��"YoXm1��y�:-�C�2)�n���Y�mkƳ;+� ���އ�Ē���vּ�Φr�>���:^yQ�j�,J�� �EA��y�5	���ȗ��Qr�}�MM�,՘��֡1MsxrȞ�Iur����]�-e��w���`���6��� d��$�q���F¥b�)z/F���`�8����jb��)�o��9~��+���ρNG8%KN�Hˉ υ�9����trY�Y
E��)P�6���DKNE��=���	���D��k�M��P��VSe8�V&y��8������[��+�-����
��x'�J�������P
������;DT��;�����p?)�C!����D��'���	E�;��g�����;��д��Q�Գ������Y�\=:�6��
:�ۘ9W�~=t��g�����9��z�]@C��I��z1a^1萃Dg�RM1�ع\��g�����4�]���\����� 7�r����%_���qRnl��N��j����AO�zpmSg�:s>���<`�=6��t��;���_��Q0��][%I!�>v�}�
endstream
endobj
8 0 obj
<<
/F1 10 0 R
>>
endobj
9 0 obj
<<
/Length 359
/Filter /FlateDecode
>>
stream
x����j�0E��
��P��P
Ml���@�E����;�S��ID��ca�cX2�݇��g�lIdR������Ƽ�_�ڿv���f�8�b�'s;�!���</Ի�]� ����޺a�v�0
6.�\@BO ��Q��LE�[^ �u#�( ��%ɴEF�-aus¢�uX��,��Ro$�=�*�'*�k���G��s�.J��]���Ad_Zob�����g����j�eW�4�t=Ӑ���4j�u��ܵح�>Xw�>���\��M�q��n4����KE}�j�VӔ�#���>5x�i�ژ���;5��T9����m�j����G9����?O��v�C��f
endstream
endobj
10 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 65
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600]
/FontDescriptor 11 0 R
/ToUnicode 12 0 R
>>
endobj
11 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 13 0 R
>>
endobj
12 0 obj
<<
/Length 502
/Filter /FlateDecode
>>
stream
x�]�͎�0�=O��t1����H�d"e�5� �H By����R���|��&�v��_�o���b�����6��6�S��Cf���vIW��^�)����㶄�a8��U���n��0O�n<�OY�u�����c{����4�
�0,���kӅs��s3}i�!�Uχ.���s\���1��ڒҎ]�MM�f��lUk����Y���U%�����f��6��ۭcv��h���5W{�Y�+͵����"�0�#���y�Y6�oܿD޲�F�1k�;��칏����~��~����`����~�}�d������6��K�ǹ,��>��N��[d�K5�_U1;�=��
G�5��0���ͥ����/ap�����R�����_k�_k��蹣_ސ�_�E�ǹ$�q.I�ǻ���/�lB�����'?�.�ך�w��6���M���ߩ-���~�م~A������,K�
����8��>�qu�u1}���?L�U�����
endstream
endobj
13 0 obj
<<
/Length 10936
/Filter /FlateDecode
/Length1 16496
>>
stream
x��zy|U����޻�tHW�$��	)B҆=i�&�0����8D��
(�0���tP��qy>u�ݙ���0n��9��
��soWB�8~����������zιg����HsK�Q+b�T�8���X|� �-5K"b]#��y��g�,~���W�!�z~���ukGl߅��!���`���W�2ʂ�hx=4��:$ ��A}P��ȲD�����}�B5�Ĥ�v�GI}q`Y���E(����������aP�DH��)��Di2B�>$�M����;���:�į�6_��CQ u��xA��hu�8��d�XmvG|Bb�3y@�Kt�JMK<dhFfVvNn^�wX����u��1c�q����?���K�U�{�7
��R��/�Z���XY�-��I�:�x���}�(ݫt�G�FO��~�O�7��h:�v��hؿ{ତ�����c�P-C��{ ދ�܆YT�"h5� �e\;��<]�GѫX���̃@Ã�c������vt �
��ᾛ40ߠ��X��<�����jf24�
�����\tXXP��T�V;�CwA��o��z;�u_�7��@I��E3��X	�̺`5Ϣc�mc�\� �Ĝd�]���;����F{��^ރv�\����w���K�)H�}����oQ#���#���B�d����s8���Ԕ;���6-��Z���a��s�O�G�W�rT%��ꑍ�=ո�U�ƏA/^ �!鶹s��3�gL/�6u��I'���+)_4N*;f���F�2bxA^nNvV�����A��nW��l2�tZ�Z%��`�)FquI�M;���(��Kꋳ2K<������<�������b4�>��Q	F��4R���zGb�8�&(<b�l�G��s�WBys��/F/��Z��h%*n7̠TjŒ�oI}[I5Ј�u���AmV&j�꠨�Rt����i�\2��A�8�VZ���M�,)v�����	Q���v��dTUQ�b!m�3;�6u����}��6p{e���6���m]Ԝ�)�Y�E�<���D3�I3z�L��G�T�Gl��r<�.�o	(-B��;D�Qf|Ϩt����nk�yD_[u[���u�G4y������`7*��/ltF}��QSu=�W��1)j�>�2ʤ��� �������6��)�w����݄;$4*��镱���;�")'�e�IOgO��������N���l'�W�E��	�����@�u>h�B"�)j�����Y���?+Uj�(�L�Y}'�ސ)m&Z1|{\r�4�E�0N���Z�-�O  "0�4#�3+�R1��"�������5SaFs<MQ���W������J:E������eV4��ڕX�V]#���L�<����ۇ�������d�c<hYZI[em]�U���+���	�=�A?Q;�А�N�~�+3+'�{&M�Sy�BH����RKn�t���Fթj��q�~h��O�h�GU�j�L�p�J�h�X���g4�"���q��(O�i|i4�T��R���}�2��0CM�Z��n
:Ԡ��Ki�eQz����=�bT*�$k#�\V�Ay��jf�Zf���{*��Q_��/s���zo����	=�b��3��� �( P>!��
K��������M`�Ԡ��%�s�(�3���S^9��r�s�eA��EY��ڊ�=x��v	�/�Sy�1����G̌�.����"l��!���TDR!�f@EM�;OH��^�6�zMF�M�ӆQMk3��QDb����H=�9hS��Zi��#�2I�KjI#�8�َI�QhybTF��qv�ì����k$glD+��b�����bN�sz����KB=����(�J}[��r�h����3������,��<E������Ү��[A�eQL4`n�LRLz��f�D$���f�2�[��j�2d*�"��b���$�9�s�l�#G��fo^���6�n�{ˬ�a*s���,�m$P�S�쯙&��(���������yH^..p��T&��o�����-�� 
J�f�IP��^��&cԸ4Lo�U��f��\AX$�	���p^�Z�� h4l�_cE�f�Mȩ�cޝ�ޜ�y��k��. �,���#����&�hUec�@�z:||�����L._u ���~�9(_��l���	/��L��>��{d��5@�n*ҡx4X�Y=PB��X�טX{��u I(�0���|fB����(�m ��p��_���׫�_����m۶��¤ �sx6�x�(�]�����������tT"t���R�\)F�Z��<��Y�2��h5�.d�����^��p���Z(s�r��-f�yX�7�������؃�ƺk�8i�A��X?�r���XRw o\��ه��|��Q�����r��U�.�s����~�@�f��s�l��+�y�-Ҁ3P��4hP��Y�7ہ^��q��9��%��3��Ly���q(Ħ01j���H^�}��`���w���+/��g�}�=p�
f`�[�Gd?��yk��ӟ��ǟ~��[$%@� ���߁(�J����Iuz�(&��<���~�E�lL%�K��؝������dG�?٤���y4���j=Y�bL�����ycz��?�.x��{��i��t=�t�����H���`���%rS��ŷ���q�kه_��0��^{2/�͡]�S�sƩ%+K�!U���i����y<w�=ᙕf<��v9�l�p��3�Ϲ53f�[|t*֜�r�x"���d�l��2�@21E*,�I�n֞&�;��[�^��y������g1�ׯ=��k3�>s䴳/�ҕ��@/6Ќv��h�Ak2�Z��a�hx�ֈ�2?r�
T6�� j10��Ⱦc/vď���A�Ӳ�m̵�C;�z�j~J��Z��[',Y���t��|J#k����SD��k�}��.Y��|M���sy#»�[�5ků��.���p��k$w��~��|��uh�4��h�ժ����U~��3F��U�*��W�X��U�!��T���׏��1�vC�lw+�~vW�`fOW-���=�e��梭r%��MBn���Rǲ���5�ٕ��4�R���6�!�̯5ؑ��/r��q�����	�{o����xV��)`����1.d��^P�`U����$w���&��e��̝Oe�j�i�C���lX�]�X�+�V'N��o}e�B�¶�ĺ�@�V��C�_��K����t�ܮ#eUǕ5����jP-�tz=����:m�_�԰,�q,�4kWv���Ҍ�#p� �Y�N/�ڙ��ׇ�'��o��e�6e����1��������P�&e& '��VU�LN@e������ɤe���+�*`A��3o^���+�*�f#�op�b�c�
n=�i��G2/<vQ��o�����Li2�����O�Z��a�a���|.��!\J����赣!�� ��kw��Vf��j�`�M6t��wZ����7?��7�>����ħ����U�u��o^�9��o״555��!:��5�#?p��`��ftě���j���Y	C�^E*
~J���k��9�H�W�O�G岊�}�|r�~���$��+2m���v2{c2�O�������N�����U�&�������j4�!R`Mi����Y��<O��;?��|��o3Q����/����c�?�}��t�;�B�i ;]�^�Z�g�hR	a�J�jPN���U��lT�{TP�<��F���O�/ܷ��=���]S#;��\�|?��z��gQ�����x6���Ϫ��/6�G��c���$�C��N�8��2N4S�NJ�[bM� c6&���ɘ�Jd�ױ�1�רX{��&�쟒΂���EXh����a����}q�~��۫�Q����o����;���)W^`���w�<��s���'�@�v#�c�s�Glx��a�ۀϣ��d��I`}�d��`�g6k�~�
'���|�m�7�K��X<b,��uc��MP��mߖ��ѽ��Z�7�u�.������z{����e񟶬:9;���;͇��3�r��'l�<�~�r�4��J#�Y���d����,�����(��Y˘��6uh�а?5�5�]�r6�_�KfoOpۻ�X4G�9l���� �CV���R�)�F�$Z��K���Y�#w5��uφ3�ښ���tݪ�6��Ĝg����wm߱�����/�>f��6��W�$x��ގ����Z!�.[��y��6bs��΀����KCu�.�j5�@�9�hPaF�T��:�5���j���v�`
���&CR`~J�D�ͺY�j�C�Ӷu�����׵G_�������/��E�X���_����@�$�+�JB	j��g0XؤDN�3Z;�;%��\jU�F֠�D�|���7�B,�X��n/�:�18,� �J��7<i���t��y��l�ڷ+��w���\��#���M��?���)НA�W����P�ಂ=�Dd���.��u�h(�)�ѱII�-#��'t�&FHe�l(4�$;���>�h���i&���)7�oo��G�^�ݻ�a~P�a��ߌ���_�l�w�/}l�\���]��=-MK71T���{W�J'�]�p�ڂzc����8T,��8�G:����v�	�7@z(���q�ׁ ނ����[�\��Өߋ��s��~0��1Ysϸ��/��e���p�Am�_q��ŏ����`��AV���2�Nmb���lO�K8��6	({��3��l�� �b;s�[�w��_��)�~�cy�p��������=�nٳU�$0�g�߅�f=8����>��_�񵷁G'@�.�7{�n���Ir��vR�8�>���
QLO�`Ƌ��z��ǔ�{�cˏ>��ꚱgyt��L,�n��~�y���:���� 2�i�X���Դ��t������v<d�[��`!3�'�G.0������|)�q��\sg9���K["T��׺q�u�oh�4,�8�^�c��͘�@U���>����K��3`�^)���0q�IZ3Ĥ$��8x#&��	t�U�Nڀ`��)~^�	/�����)�s������3!^H<{8N}?�Ϯ���B�6��V��v��ʤ�:��8-���9 lp�:k�5��o�Bdi���_q�M�L��m�K"bU
��hhA�1<���[��W��x�z�ʧ�˗w�:�g�9�h�:�y�|�p'V<�h9�?��\�Z^ݼL������6�+�s��j��l:�æ����U�LQ�e�U���� qqo��9qL�6��q�&r�yŭmg�{ �W9�Y8ׁ�j�0)	<��h�,�e�:c�p1ĺ�Ȍ�ua߼��u��.L�6������z�0O:��	*+t�,a^��he%����+R�m�	d�j��ʯf�C�p�����<�DG�9�07�`w��?�/��4>s��r���O��w���%�%�"w]�Np�ȳ�b�	8;\J��!���;,�r�e~���@R����cI���yނ��*�[|��i�g=xWk���Lz���O2o�v)���s�[ ^OB�RJR	�Նl��&+FV����dm�vZK�-љRj�&$� �p����Z�ڪbUt�&a��ļGU7�5�V�	�n	J� 9�lhf���br��u�#;v�v�󩸥�-��1)�n<��0�ᵏ?=�p����~,��z�bS*�&YT��2�ZC�X�I,��������Sr	7�;xm6wp��x�W ��K���p�V��0l��YnR7�l���9⇏ m{�uY�&�\�3��7���+f����>E�R|@�T���4X�g�r.ޡg,�L�`������\��z�bA<o�!3�K��yoˍ��7��4ڄ m��K��˧�g���o��w�q�և�®������LR����s��Vr�J�,px�xI�W�sP�i�M�&��`Q�X�M�r01F`�:r�`��pf�`�!��Y,ه�b̫T�ʯb����j�����cǫ�ǻn?����-�t}Η����E`Gv�&YQ2o0�9��=�D�m�8���.H�_:�ML� �<����������F�<+<�qs���^��֯ݵn93P�B��#�^?� wI������3�������z/��oo0�3#�dtUN_���qj�X`auHWQC�t�WuRd��[��5<���x����ڷ{�pq4/����E9kʕ���T/p�Z�s{���s1�����~��pDju��/�����ةӵ���ҵL~�C��&J�~�c@��d�ee�'��b���D��T�%�L`���S�X�obH�#��� ;��>1�h��0�)W/��<b��莽O�[xo�f����g�L�v��e���%WT��掷q]�ꖕ;�[<�E��yqg���h��<���=�����f2ȆG.� z��A�32�E�L�d̗N3� *��t�xQGs\;90������_ñ�*?Y�Ϝ��3�X��4g�����#�\�?��M�-��Gzl'sP>"��ux6��}B>�ػ.���qBL��T��D�+�N��ڵ��$����k)1�\�_�OH`��*�N���0�2E `y(���&qE�#��� �@"��#��|����5��9���=�(�(ޞ-�����x.�%��/��t}:T�e��_���R�nƃ�J��2�x`ڠT��U6�l&�em6V�1��F=6�z�Fźo��7r���#�7%a�c�3v�{��=�bХ�~xQ��qa���:�w4�����3q�G�j>����x�����:,���ܪKoo�7~�ߜ9@�����OJ��qlB�yl0"Nυ�jިw�s�!=��c� ��
�q��N��v)��5��|�����?O��d=���q�&v���[��]���� O��5�Tɬ��L�դbY���w�f"AC"`���1_\���閇]s
�]������?sf���>������)#���
���JHT�U�$�`Щ!�5Zt-�{u������h�m���c���{�@�66��^��>|��$���2P`:�ud���?:ϝn]��1^;g0����Ʈ�CL�����}��yvâ�9U��*j�����J�����0���]�s*5���#+pX�Y�`�@$���k �ƃ-hȱ����L�rV��?9+����O�)g�bw��*d�t�ʼ̬��� ���o:rr��h�*�q,�	<ϰ�N��r�ac�A��Ƚ
b�y-���˧�^�{���L<�M9��'�b&�1�s�]W��'��,�/�}vBɨ��8v���E�S9��s�n��{����/$H�C��:�z��S���|I.�x�)����<���-�-=�uZ-����|���3��Z�&&�배-Otv�v��k���gl�_��.�������ɔw�sw#�Z� ,,D:�ƨ�X��FH��7H=�}A�L�H~o���.o_������	�m��|9ğ�`�䜮]�s��yiP���b1�0X���c!�1by���7��#{T�[�I�	���`�*vr�,�l����g#���`�јJ�L,�b�;�=s9Ze��%�.��-&�͗A\��f/ҽ}�t+�U������\�����p|�IG)$���sq��M�+�[+��w1d��:ď(p��k%��a?�>����ܹSF;w���z���3Rrq���R<ðF�c\�Bh���^J�y���F�����?#
4� �9ןd?�!	��8�����#�c�B!$�X��X#��@���M� ^��
�d�0��������?D��{v
�z�/iX@O�[%�����Û������ɻ[r�7 UJY�	V��fS� �T��-1�ٜNS��ݞ��N�_�%���f�4=�wʪD�6zВ>����Cb>��Aܤ%����o�ߍ�����'��0�ú�����k����Ç��w����d�`��~y�����Vv��FVGǸb��}c���z���}M�ͽǓ�g�{�̉�F����N|��=1w��S�t'Z�j�s��"�����}�NAy'jF+�6�����)hiC'���<�����G- a2��a�+ �-\��ATV�w���m���e�v����/�p�� 4�{���ḍ�"f=e��u�>�.�k�s_�_�2�e�[�l�"U��Qg�}���4�f�f��]m��Rۦ�L��n�n���~�>��]�>.�����k��14�n�d<l�hJ6M5՛^S8T��w���P�!�kM#�)�����zy��jX��BA��Bn�H)s0�>��#z@)P~L)��
Ԯ���>&V� �e����l�R֡d�������'J9�Z�l@Il!���@�0�W������2p�̢a\�R�`LP)�(��G)Pޫ�U�*��RV�����A��������V)��-��V�zt�Ƭ���B�b�l@�4,nX�iX�k��XjZ�ܰ�>"�"���劷�B���Ps �j�֎�yX�8@�"��ƚ��󃱱�PchFpAˢ@�pM��6�,f�7��:+�&�����l�Λ�6�ŀi��%���!64�#�fhlh+�˳Ų@$�����މ���j���&�	��P��\����m�!��ٽ��aEy$�$(N	D"�p��(\@��PK��1�).�o����bm0ܰ���/���7 �il-�K`Zs��9�oh\ ��a1ln�S@���@��}q0��PX�h9�mqL�rZ��'���ҩ����{��cņ�M͡%�ЬpMs0������" �>����j-��)ИU��j
��o�|c �ci8�hI0LG7��a"�ZX�"���B�"K�5�����>tׅ#05$jka���PM�b",�u���@Ms��" eq8�>i���t���"�O6@������"�fe�ɠ�D~-T�d�&�Ӛ�?> NTd�=ꙗ��� 664E���E١�9�|�Q1j �� �N�"� �P����	-�OF�C��C�x�\���n�Q!�_�E4��0��n5�l�����Ci�BE)��	�	0� L�y�/\M���� 6�E�یơ0�	BO-�!�,�~�/�΢=���|�(�ٰI���_�� �D���!T.���
�B�Y�'D�rCO��j)T�F��Qet&�B�bk��f��i����P������.� ��\��s!�RPK���-����?�唺%��N�a�W������*�Fh'�X
�����<����5*��Ή��KT��4R�-Q(]�`#\���0��8D(�EJ-�H�MT��k*���Co�����E�]�X�b�Q�|Ş�R��]?���Tx.u���ϛ��)K���tM78�E�D��T�R�Z�|�����UO�$@�T����p�VY%��D[� l�8�(\�a6���?1ƽ�ZJ$������R[K�B��&�)�b+^D}үz�TG5/��Z
-����&�`Q�j��{L�B0��J1fY1������!e^�M����R�6�Q^� u�M�����(֓�М�=���D9��J�{iY4NV�@c������I��7�L=G��?>�s�M����=� _�M��ic�#��0�e6]��&�bi��=��~�3.�C^8U��s��lȅ+���4�l�O�'�������G��V��gv�Յ�e�a�C�l��R�����Xk�˅V#�1\��h�'�^�ppiI���bTс���!���P��i� r� �@<��z!��J*P��l���`�?|C]_�
\[/�|�2���
s�
�w��T]	]a�E�"����v��4�W_�q}�E�����g>��3,}�s��|��:}����γ�y�p�y_��$����x��~[qn̟*>�Ig���\vX��cX���� �c�T�v���?�?)�����'������z5��W�ӯ����\M��x*�T�)��T�)�x�u��9Yx2t���s'�Ϥ�Ď܎��������L��c�x������\��1��\�sW�c;p��q����e����Q6�H�f�3�g��g�}��9\x���4�<��!f\6�|l�u ����ba&Ɏ��T�i��>�`��7�4W�.i4<��#�Gh�<h0��9ڵo���Ѡc�)O.�׺pv��;��<���v��I;N��>㎜�;V��7���(����lߜ溿��un�݆]�r�1�m��1h�i�����q�&$��-�[�i��6�6����q�kS�&V�d��L��V�C�p�ݝXw4^�� ��d�m\���0q�k��1�ukG�����{/6���es����`i�F��|B�\�p%ᄊDoB���V �j諂�D�y�:�J�т�&��S�ݗ��9��[*x�Vp�,h���s����8'-pI�����Z) �(s��L��H�n�I�S��)��&�ɾ�I�RWYvJ��D�� ����:���|W|L��c{�#�^a��
S���K�`_��Z��Xh�2�2rFc�q�1d�j<g�6�
�튑!px��ok�Y��1�C�=cRTS67��GS��]�>'*����9s+�1��w�fT4`R4��2Z=�?)Z�Z�`��@E�p$iɈ}�R���H��B{�B=L*8#�����HF�g��=�X( @���MaR$#�a��"Ha6� :-�� �p�#L�w�����K������������y
endstream
endobj
xref
0 14
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000392 00000 n
0000000115 00000 n
0000000549 00000 n
0000000604 00000 n
0000000761 00000 n
0000001879 00000 n
0000001911 00000 n
0000002344 00000 n
0000002771 00000 n
0000002971 00000 n
0000003548 00000 n
trailer
<<
/Size 14
/Root 1 0 R
/Info 4 0 R
/ID [<D0525B4A0BA8D19012B375531A432F4F> <D0525B4A0BA8D19012B375531A432F4F>]
>>
startxref
14576
%%EOF
