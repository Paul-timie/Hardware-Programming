%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20220929002115Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R]
/Count 1
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 6 0 R
>>
endobj
5 0 obj
<<
/Font 7 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Length 874
/Filter /FlateDecode
>>
stream
x��Wˮ�0��+�f�aǶ����#U�xH,��~�3vU�:	����&��3�3.��}?}먣�$vs�w!�ϗ��������^>����}�}����wL������z{�rZϧwU���C�%!%G�
)�H҄!�Kf����+��hHRq{S��?pb����U�/w���ʎ=y�y<h�}Ěp/<��4��8��l��p]xA}1݄�kn"�+oR<���	OY���V�=���� 4"���]��Qlv a�yot@��  6�f�p�q��Cv*�"�:���Vj9������{�D�� 5�k<�#���������
G��"�,��ɇTw��i��v*����&֪+;�ۙ�"�~۸�6�9�k5n#�e��kւ��E�|�'Y�����
�~�\r1޻�P.brnm���B�K��B�K�6]Ȭ,�Q*���\%�2GN(�Q�MیwuS��� P&�L;��Ӑ��Rw^ZJ�S�?�,,�����`g�����@�L�g]4=-ތ��L����ˀ�J����ɟ�'?Gˡ���hRS�)�>E��g��Jz.){.9����w�c�xf{[bY�q�,M�>k.�"ј@�5kW0s6ʌ��+�)����;�ɶMǡ&��^#�lH��ͧ����-�̘����G�,�2[!��6y�1/�4-NO,K�:�ݳ�r�qܬ\4喘Ԟ��ȓ�%��I�&����]Ә؁d�gR�M.�j�lqq6u< �q7誤Ѐ��='�n(9.��sJ�$�Ӕ�S�����	zJ�r=�#1�u�Y9q��y<�Q��~\��inԸ�}��u)��!k�͚tm{�+b��el�B��;�����Bs���}�D
endstream
endobj
7 0 obj
<<
/F1 8 0 R
>>
endobj
8 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 62
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600]
/FontDescriptor 9 0 R
/ToUnicode 10 0 R
>>
endobj
9 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 11 0 R
>>
endobj
10 0 obj
<<
/Length 492
/Filter /FlateDecode
>>
stream
x�]�ˎ�@E���^N#�������"���!��m5f�ߧo�N"e:Ʒʧ�T�=�������b��������/ØYg��[ҕ~w�v��X{|�=��i������m	�駓���_C��0^�ӏ�1^����_���"[�M�ϱ��v��^}�Uχ>���s,��x��8��T�����/>[�ڬ��u����{�c����lC��-
�[Gv�,ʥ�K�z�Ț���7�݂_���Wf^�eـ�ؿo�o�;���ɚٳ��lr	��L������������h����K����O�R3�s��o0+K�g��_k�?���_o��o���_�ӥ��ӥ�k����+�ץ�c�.�>���+�������쒿f��f�_b�Byӿ³��%�%�g��x�B�
s��x�п��+�W�����!��B���_�^��q4X���J`g�����!�5�����f�����4�J?�H���
endstream
endobj
11 0 obj
<<
/Length 10786
/Filter /FlateDecode
/Length1 16236
>>
stream
x��zy|TE�p��zM��Y:�o�d��i�@.!ih�4�I�tHH�t��@ª"���
�tPApy�8���3�=a�faEGr�NU߄�q�~�����u��:��:u�:�:Ѷ%!�G�ER��`+�ه>���Q����|!�����92�*B�6�T/.X��qn������7��o�Q��P��Mа����P�	�C�G�r�5�>�����Ŗ5?@�ER_��u)��E(��-�š�% ��DH��5��D2B��'��m��Kۿ�����І�K>z RgX�Tj�V�O0Mf��fw$&%�8S��D�`ϐ�̬�òsr��
��ËG��e��[ǌ���������|9��:���F#Z�P�R��S��Y���T��ŋ�Ut �Eot�ҵ�=�N~�BϢM�څ6����Q���B�Q�_?���.�������Eu(�V�.X��uroȕ�<>���t7�fv ;���q���3�g�>�]���=��C-̓l9� ;�c*��X{*z�Aw��5���2�Ih��%�{�5�;���*P�mJ�ѝh��tf�J�f��y�D�6������1F��0��S�ۀ�j�=#7ɻ�.\���6�����|93�{.��jA�h>��{n*��F��i=_3א�s ��;���a� S�`Ц�z��ur�1r�I�0�Z�j��\�q���;y��cЋ��oH�m��@M�̪��ӦN��<ib�m��	�㥒qc��:z�-#G����def��v��lf�ѐ��j�*��X�1���cl�h�=�`En�X��T��S����Ġ����TT�&O0&։�(����b�l�i�)���&qC����3e�Ϟ^��2O@�]��
s�� �fP��by̷����hĝ:�τ�67uju � �eyZ;q�8L&�|t'��	dY�iy�!�^S^�t��9cO�B(ʘ0!��(�fB:�(v����eB������ܚ��lyGǺ�9;6�S��$�y(��)+�e��g��3�ƒ8Ƨ�<bǷ��xa`KPi�M�"Ƙ	1<��M>N���}u�����������;Zˁ��_(�z^���6b��&<:�l�7cr�:}NM�I��MAh�������7�����v�	6vIh>Tb��k�u�wFR~v �ԑ���=�j�����7����\U���'6xʁ������]�`<���;���a1���t�TMlhc|0	f�� zC�t�h��]���2�q��<��:�oiS ���qE�Y�� �����;�aF��\F�����l��>��ʛ�j�eZ�6!���Y��rjWbyG]Y���3��(����.:_��#����	�e�5�1W���Q�q�cR $�ԄD�CC�9�r��̬�\�<}v�-
!���K/�	���G
S�����`�	D ��1������ᴕ(n��;Q�h #6T,�)�H} R��ӄ�^l��	Nw����0�-*�5ajEo�)�P�~N��M��ID��O��4�1�_C�F�C��0��\����~�6!7t�V3c�lg��n���j�M�{���grUA�Q"�|b�n1;�/ ��+����AwtJ1���gbC���f����d-��'�,���V����wJx}�욣&���Ϭ9�`fB]i�s���Р�i%��"�
�4*j:�yT� ��r����0�m��6�께x�)�P]HB�p��w4m�x[;m��NDX&iyI-i$=��8;1i:-/C����=N��N�5�6w��N�䌏h�R����7���]��4���J��%�	��J��@ee���.@�9@4��c�3������*��<��������Ү���A��&0��&)��rv�.I��t����V�����Y�
�Iz�XĪ5<	����1[�Qf��[X�5�ͬ��^�2�e��\�0�e	��T�>���$Kz�;F/�1�(^6ERX���v<�)����K"�;{.pK��ȁBR��dT�$��'&!���5.��l����!�@�	~a��	WA�
�F��4VT�mFޤ��;��Y���F �#뚽x����-12�q��lr�VU�f��gc�'F�yH>,� �$�UϤ�j��O2��������7ᅸ��;�߹V&�_�O�"JDY��"葀��5F@cb�� � �PRIv?b�	vx�g�`�9�$nⵋ�G�_�^zu�û�m۶g�K��C�'�d�o�W��~��ǿ'Z����ʥ���LPJ�+ͨVk�4YC=���RF�Ioti s()**)�z��C}���B�SX�6�i1{��3��v�8�-r$���f���i���fp�ԚYV&+\�����S�����ݏ�U�[U�8��a�샿��'��<ӽBm�<�+���1�E�f���I�;���U;�?�1�</�Нݏd�C��L�C!6��S;����]�U��K�!��\Ѯ�����+��ﾇ�]��~�K����#8o}Rs-p���^��ӏ�z���d��;�it�19Ţ���#[Phɚ�X����p�����=ɼ�MNNMu��&����� ϫ�d��q-P���Ov�Hw��Ez�H�����1�Bf��G���2-n"�#�h�U��MIq���0G�w�yt/~�����&�<���Sú��n���KW�ªVSs��w�y<w����3�J���.�}d�~ƌb�/�N%Þ�P��H��4�l�m6P&H&�H%%7)��ړ�$zGP�a�#+��(�T�a�������{^�ս���3jڙW^�·�KA/6Ќv��h�Ak2�Z��a�hx�ֈx 9�*��)�Z�,&�/�؋�#�m�xȤ���i,�X=G5�8.�8!�ҭ��.��q.���\{��q"{|^-�fJV��!_Өyn�ވ�9���Z�+n ��_9�<Ζ?b��M�"�|���͒F�b�Zb�	��6���y����_����*���O�� d��� ���4*��n���n������bvw7��/�-�~D��i.�*�pi�d���.es,�e��Ѹ̮�B�і�$�L�@k�#�? r�q��E��	��^}���zV�ݑi`��b��q.d���^P�`U���ϜN�2�9�{�����:���;��e�ܳ�k7��.
V���5��'OǷ��`!f�Xsb]s0m�~ā�o}�%��k<qv�!�e�������H.�^�5���N[�!5lKmD*�ڕ�d�4���,~�3��v�x��a�)�5���ooٲ�M���ɓ�5�_����4M�IB(AP%[��֙�����$���ɤe����e�i� h�wȟ7��l�˕r�z���78j1�1x7�K۴`Wʣ9�� �p���r�}�y�"��?�L�]y����.�3�l���ø�����;�kGC%�A�#��H4X�̌�դ3
���l���L/9oQ"gomx����f����{j��֯_�9���w�;Z[��������τ5GHN��f3:�z��5���,���!f�"e}J���k��9�H�W��}�����}��j�>���"��;:�r���ۙ=q�zQ���L�j����b�j�����cg5��)���ll�s!�ps�'�	'?��|߇�21�%y_.�_��_�k�E
Z	z1b8�L)/%Yo�G	���Iؘ�Jb�$c�+�����j4�H@�b� �|�ͧ����v-4��&�p���,�Ag�i?|���K�燋G6�{�����.לg���w�z<�ó����`�� �c�s�lx��_����yP�t�JY������H@o4��{�����=FA���ݞ	�U�&hU�������?o�6�
���7�jI�x����8�����O�:����G�c�^������|s�5;v�W��ʜ����m�����f/F=g>���=v���[��Mu�� ���TI'l���dp%%����F[|��{6��?Ÿ�n��H�2(,ܐ��l���fm$`V���óק����
�u�8<r�=��ѕMP��m�V���=�:��6't�.��ѥ_�|w���ݒ�ܲ�ج�]?��|��'c�/�zb����Q�t9Q*B�QI�\mfB�}pBB�`�]��H��Y˘�$�6}X��H =�5�]�r��_ԍfoo ݷ�x�HFl�ν8�Cv���V�i���Dk����ß?�y�����w�n8���uͮO׭�{C�J�yvo^�k�n�+�~��˫_�s��[��	<��yg��߆�lk	����Z��m��"�� ��`�M&���z�a�&�	�j8 p��p������ܼ�y����$�W�H�|���X5�)���ݾ��Z��ԏ�~W(v1G*2��	z�.�<$��ad3�-k��9"��Y���}��^b	7lb^?W���j�X�2v�+*�NV�Y�͇d���K������Ñ�9���I�L~��v���8 !�\�R�����ksj/��m�e�y����_��y�2�|���5�� Ǥ��ԼQ�����zNS� `�%����'��N	w1خ�nv���m�ݿ>&o���*.�#�d����-��Ʉ�p���P%�1,�L��j�9�hPaF���ӳ�x��p�$**qΛ��k7��{�!��t�nփ�l� qڎ�3����o�w��w���ÿ�����|�{)�C9���m~5�5�JB�ÁP�Ze5%$�$6%���֮����`����#kPH��P[�;�o�%XP�6#�
|�Z�%6v?�J�'6<e���xԞ��s�Olú҆w��I�?�w}7�1�Ňgo���+q�}1]�*S	.+�1(Y.3˥w��A5���0:6%�ab�~b4�����%����DpW�C����>�f̠�.��pC���p��|'6���o���T샔}���}[5w��[g��G���}ڳҴ���U>u�*[Ť�c*���KP_�<x��ʤ��H���z�6a��f����U�%j�
�x���WB^rZ�gL�C/��[��������r�[xp���|��-�ְu������K�s���hiP�0F��b��Z�tj��d{s�xb�?��Q���$�̈́f[��������p��w����/d�������e�=�i�C��z����$f���w�ǯY��0F��O������� k�%ɽ�NJҤ8�v;�vG�]��?��as��(�7�4����z�KJ�6��凟�Fw�ؽ<���\.�����<����p�u ����#d�H�1/J�����$V6;�������,o�s�����p�}�ӛ�[8�/�>n̖k�\�US{qK4.�; �b؛�D�j�F���"������	*-�9pEl<�&���2-���r�`���:��O�'�W_�{�ȯqvJ��'�1���a��d���`�k=C������]Ұ<�0z%�!�3c�TU����?���?�Q]m��jGi�/e�⬬N'瀰�%�)֔ڀ�
���F���#�G�b���@�!BƤJ�x8=�A
��~�|骜�w�+�V>}D��s��?��cױ�Гx�o��8��d�a�����u�궻���)����gCR"�X�6�Φ�;lZ���p*"�P\�޺���� ��q�u���K��o���h�ϟ�W��qF^۝ߛ�Ú��:���R���F�2ZF��0�j�A.��=n�%��z��|7va��3��H��֛�{2����Tܵd)�z_�_K�l+YI�L�� ��ƛ@��VkjV 9�O������M��"N5���]����>�O_��I��;��g�Ο���-���.w_|���D�Ŗ_M��R�����v��\� ���YI�r�10� ��q�[�T%�d�ν7��w�w�����N}����,c�3��bzy�s)�IJK@�[m��Lm�bd5Y묭�v�I��a�y%:�*�֤$$�r �T�T[U�J�8L�p�w��*��F��j����(P�;�Q!�@k0s�?.��4�/}���h��x²7�ۃ�4l��m7�i~��O�,\���U +�u�bS*�!YTs�!�s�zp\bq�6 �pۙ�<.�sù��fq�w�&� ��^�1M���*
�huz�k���r��Qe+R�͑8b$h۩�d�),���r�S|�������>E�V|@�T�4X�g�r.ѡg,�L�`������\��z�bA<o�!+���-7n��ވN�L������\:�?���W~��}/�/_�I[fJ�_��_{��)�ϲg������<�����%-K�Dz/��<��`�+��
xō��iP�����0�Ց;)#��k1k�cV�b�>�c^�B���7/�Wۍ+"5���f�x5�D�����~��h��|�nz?�\
vdGnѧ�C��<�cK��6S��Y�8�S�à����'~�Q�5�z�7�^�ͨ��9n�7x��w�}h�=;�-g�_�_u4�G��.ʁ�s��>}��ǟ�����u���~f��*�����k4�N�R,��j!Z�
���b@ʅ�bz�)���\?���o�}�{7�@�-p��kQ�"�� �������9j~�����?;;{��$��Z� �����F>���v��{!��4�w�39h��%���R��:x.7o�>�M��%s��6 	~��ڗ�{��M��yD�^B��F�/v�4&1���o~�GN:�{pϓ��[�؆þ���s9ǒ��\��x���+j�2q[׻�1}���m��[<�a��-��{e{���h��B���3����"Ȧd�#�d =�� ����"rgJ���'�������h��5vrGd�75�D��6��Xkm���G���D��&8����(����b��X}J~G~�ч�����q#����h��0������ȩP��a��(�
C����v-�&ũ��"%'�+�kII�Z�P���c��+{-H)I\�.�	u�3J�D�#F'�M����X�gG�����1\]�@��1>{��8�'�9�v��[�|]�s���D���nZ��0�tɬ��-�դbY�V�C4�.���h������X��ck����~scv���N�y�C�G��As�Ӑ�y�h?�$$�h�� ��<��Hb���4T	E���2�AN��A8�k�xzXڑ�����<{��L����3������y�-T&vX���ݳ�<�,F+�:�rV���V%��)���S%'C�h�����1:��1c��2�<�g�ľk尙$/�Z-�#�$1>����魣2��͑��ܙ�u���p҄b��l���@��ߏ�;?#�j^�6���d���=��O��$�Yi8�h8	�<�Rs�=Ұ�՜EFRDZG��!q�Nݡ�'\3�x�y
���!o<�?���a�ܽ������s�=�v���ف���Z��c���F-�ʕ[��L�DO���!��<~��'�8~� c�/�e.�W =2�#W.�(~?�_ҋ_�ղxbD�?�����b61�^��]��ɓo>�̛'�����ȷ]�;~'`=~��W�Jʿ�����,�R85�aU�J�S)Q	ihm����^��䏄(�ͭ��[ԝȾ~�]6��Kٽ��gt�(z��� ӹU9�HP�1�8�/��*�$��B`�fP�<��d��{�[���5�e?��;��������|��4.��n{��!�K�rX���.`���Vnw��SXN�8* �y.P����b��v��c�2�C>�)(~�g  �	�`�9[�}���o�>�Na~O�]!�b�=ȭ��Wbz��<��\E�BG�,�vV�q̷�+�?�oOX�t��)�\�gq��}���'��~�߿:���sg�*<�;�T�^@��B|�m���kt��h3jC۠��$�dh5z�;�Qȁ���Q�l��%��b�}��u���C��j���x;�o�~Ц(H�;�4���n�?x�`8��Y�Ę�l#����+�ڸ������
w;Y%�6�>U����j�RM�旚���>�9]��I���k�V���R��^NhL�'�-C�a�a��1�8׸�x�x�T`�D9R��p��1�|4�ڣ�$Dz�pK�n��!���vf@�B
�BޱH�9s��ȀR`��X�V�NV#ĤqX��D��p�LQ`JeN��gx�'�bV����9���(�-3��y�EùB�`LH�y�ʭU`�=
�BW�WX���C
�A��X�|���:t���X��j�
��j+�����yAs�yE�AlF�b}�uy[󂦨�U?T,*(,o�,
��m��`�9ܒ��p�"q��Fsĉ-�y���C��pKxFh��E����PKC�M�opS��P[��Eyy��7m��A1�l-��L7$Bl-h�DCm���"V�U��`4��-�̾����C��>���p�	�\���9��\OV����ߏU��Ґ8%��"��`��&��D�[B9Ⲧ��&qY0"6�"�Z�{�rq�,z������R@�����B���b$�#���F�m
F����m���E�������� �e��&�~[3P:5��@^/5��F`�ؼ��-����o�Z`�`Cp~��(�j
��m����epCl��/i����Y�U���Y	/Z���-�PC�����&��៑-5�ۀ̆hSn?��-Q���w`X�~�b",�u���`}[�Z��eq$�)m���lٲ��"�zO`������֐"�6�e�JЁ"�%T�dU+�i��'*r�^�,�+T� 66�F#y��Ey���|��5��n��'��O�A��Q�����ɨ&hQ����BxDt�
C�"�/�	 ��,�R�aԂ���O�?b+h�BE���D�_*a�|��WDSh���1�z��x�9!�i�3D��Oc����iO���(*�o?6�6&��8J{��)�?��0�?�	ƅ��"�����ஆUt���$\���Z訙?��4X���S������.�1�nR��x�F)h��z������?�U���t�)���#���e_q�K�Z���cPC�n�p��b ֢̞:'��Z�27�Ȧ�Jn�B�Re5��F���u[`� ݵH�%i��
�r-He��b�ұ�о��k[<��:_��e�:���Of�y:�e��T�yנFEcɪo����R)���(�
R�3�u�t5Q=	R)��G)��\kPvI�n�-��-�k�R�d�Y�+*c�{���Hf�7�w������8MF-RV��x�I?�R#ռ87(����Fʛ��j�R� ߸����K�����p.H�V�R�UhYL-���a+�e>PG�yT��O�b=y
�����]����������@c��Z��oI?K�Dx�J�9Z��)�o�@l�f�Y�޴��66C=J�P^��=,��i�Be<�����G>�3p�SSP5�����Ȇ\�J�Ӑ��j\	%����1P��񣡼�,������<<��a�=^T���ն��o-�y�j�7�'ޚ�P"�u�@�o�B�w��.�{x,)r^@=���f\�3L �P�*����T�n��?���/��w�0�_�k�=�]b×�^fN\�{/c������,� ]`��}=�?���ꋱ�/�Hs���>���2~���|ן��\'νw��9V:��;�Kr�64�jl��c��c�X���O��xv E����ö���ȅ�f���q�R-~������'������}#�ƪ7��������X<^p��q��x�q�x�u��?Vr,|�б�����e�Į�.WkW{O~�I����`��H�������K��.��v�)�@��=�-��b'c����C%����ŞcN>��sL����̞g���`�'`#*����	va��ؿ�nw�n���_�2\;�����G��Т�a0��>Ƶw���1�c�)��KY���=.��C�Olg��
}�v�^z���`��%�z���e�Ga��D�����z\g��mص-޶j�����[Y��֤T���`3ms���f�`6nrm���J�LV��$�"<�='��p��;J �o��6��pm�4Ƶ~�X׺{Ƹ����s/6�#�Sp[��Z��5�/�	�r��������I�*/[-�d렯��=��+�G�eM��1��5�W��l(�E�j��\��~�9�ed�Q�����.(�|]X+��~������4���4==�����ĕ�A�ɾ
��;��x�c"V�m��᳾�>�݇���Qd�6cc���X̀�a��Tg��e,1�W9�1�8�6n5�5�U%�v�Ȇ8	�ׁy܅�uά�Ξܥ�19��ω����*�ώ	�c�z���N���ݼ��+����
L�5  � ӠN*D�����+`egG�P�
�e�~0���H4QZ`Ԣ�K�;;�H��`@o
����0�,
�q�ix�.	��d�;"�zL�8-}���S�]�~��_J���
endstream
endobj
xref
0 12
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000386 00000 n
0000000115 00000 n
0000000543 00000 n
0000000598 00000 n
0000001546 00000 n
0000001577 00000 n
0000001990 00000 n
0000002189 00000 n
0000002756 00000 n
trailer
<<
/Size 12
/Root 1 0 R
/Info 4 0 R
/ID [<04F0613814EEEA8971A03D299B21C90D> <04F0613814EEEA8971A03D299B21C90D>]
>>
startxref
13634
%%EOF
