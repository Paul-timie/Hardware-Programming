%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20220929002114Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R 6 0 R]
/Count 2
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 7 0 R
>>
endobj
5 0 obj
<<
/Font 8 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 9 0 R
>>
endobj
7 0 obj
<<
/Length 1033
/Filter /FlateDecode
>>
stream
x��XɎ�6��+t�AS)�@@��� �Y�d.������IQ�A�-�fիW+�Zn����PC-I�t�m܄������ן���_`}��2�.�k�&H����[�iᆩ���3��_����̷��I�ۮ`���#O�)�@RC����ǯ4a���3A]�"��C=����Zvaޞ����{��.���������wxy��T6�fa��_��_UW��{I�@�'�yI�܉���~%J�8
�����KU�e�8Ⱃ⌲��k��*��1'q �0JH$�	W&BhY�-�ߎ�'D����mbX'�5	<GR6�v�Gj�$�C&ہfz�'b٨ꡮL�zh���Y�M��X���\����]
��T婪��V��bw������'�U��zE�%􃯚I��M��X�Ԉ {Ai�R�

�<�E��U����3��$�:�W<_媞������u1a�s �F(� �����4���|��P,�B*�{`	Mj�a��8Y���7�*���T���ߕA���;Q�Z
���'#_ZMz��h��*4�Re�]�W�4ʰ�guٓΡx���s��x��i�ŉ�4�r��� �>U,Ҙ �f���� �ܕԬ�X��\[u��]�|g��f,��P'^�/���;A�d|��\�R��1�r��K�|����x7�L�xT��W�����?�O}d�/��V��8�9S�XX@g���T��*1kpr�4�'�Z�Y3<��A�:-R��6���`��`���m ����
%���s^t�ᄓk�w�S�inWU?�q��/!�Zgr�ӼT�{�IO��fj�&<��9���4���\�����(��}�Vf�Ç�n���1�R6`��P���c��(�8ꡛ�����Dd�_�6��c���_J�̯I��U���0��#�~|Ұ��*8��I��o��U�����6$G׎E>�UJY��U���u���I��T��m��5�����1��|�Eڞ꺲C������?�;�]
endstream
endobj
8 0 obj
<<
/F1 10 0 R
>>
endobj
9 0 obj
<<
/Length 647
/Filter /FlateDecode
>>
stream
x��Wˮ�0��^wA��RU	��_)R���+�n�� �`���jb;6s|�x<����5�W�n*���o?�o���<C��W՝+ck�ٺQ����
A�~�3�K��O~l3�Gd"dfM����KSfr�{���#������w���.(4�-���� ��,�5%`y��!��<�4�WچR�g�y���2�$:'��p��� �N��pA��`7�Y��ܞi-����cl�Ȍ��-n��~�7�1P��y�~)�#���˳ �?�%9��G�n����2�󠴻���i<�مl%m</=�)b��V�(í��h�{�̳.�0�� �����Rt�Y��3�P��	�=����>L4�'�Z��%��G1�4P��Xh�c(����Gl<��@��O�M������aܜ����3�m����qJ7;ϻӦ�4Eb�L+��,K�@�S�De%B�!.�싘�
+���v�H�r�M����e,G��x�7l�e�z�	��ȶ�{��N�=+�)%MZ���Y�%k�c�� �eF�5eEt�����Z�ވ1:U��0�E����aɺbL$W���1���~հrn�T/��c���C'��&�,����H�'j�>7/{Q� �{��
endstream
endobj
10 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 66
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600]
/FontDescriptor 11 0 R
/ToUnicode 12 0 R
>>
endobj
11 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 13 0 R
>>
endobj
12 0 obj
<<
/Length 505
/Filter /FlateDecode
>>
stream
x�]�͎�0��<�����k`F�"e���E�L���"5�Y���s��J]}����	�|{��~ɿ�c{�9�C7��x��`N���u���%���^�)����㶄�a8��U���n��0O�n<�OY�u�����c{���}�~�kSd���9���L_�k�u�󡋗�����+�xL�8][��cnSӆ�.![�ڬ��u��kU�-�s���c���E�v�Ȏ\�E��+W{pI��J�����-���~e�+x�,����-�k�����d�ٳ��l���+�_�c�/�c���o�/ڇ����h�|,�K�I�g�����������}�_��ҿ�Fv����%=O��.�O�򇧣]��_!O�򇏣	����������������֧����y
��L���䏜%�+��#OI���$e��Z����e�;e��ޗ�N��_"��C�B�����_��O����&#��3����sK��<b�!��VL�]��e�
endstream
endobj
13 0 obj
<<
/Length 11338
/Filter /FlateDecode
/Length1 16984
>>
stream
x��{y|U�轵��޻�����	IHR��$@ D� $M�!a ��*J ��0#�+��" �9����3��d�q��uRy�ޮ��q|����^u����ܳ�۝p�� ң�"�f���� ��"�-5�b]#��E��W�f�{��}7�6!�zu���u����!}!B�����ݷ
2�~�R�;�
P��~�������1A}��`��#k^�M������q���.6��������nqS0��Re�F#�Ḿ�������y��%І�C.=RgX�Tj�V��1Mf��fw���'$&�Iv����~)�i��dd������7d�]Æ�=b�|it������gу|��j��uqÑ-D�����UѲ<U���u��*z�E�лPzD�Z�Bϣ����@���h:����h�\�(����6������hz஄�^G3q+fQ5
��`�qm�[r)�����=�3�-���)���'�����%�+x��v��|�gF�F�y���V3����������Lа�A���Z��8�
= ��={��ڐ��`�mL��h:��td@K�z�	�y�mk��
{�&���؆��x�ԢZ��D/�����"�I����h	_ČG�Ϋ��o}�Q)����o���
~g��Vr�7�Md�H+���\�td��Ҵ��\-��#�����o�ŨJX��#���?��`���\�tC�=ӧ�*+��O�T6q��Ғqc����)-�9�����:$oPNv�����Ԕ~�.g��l2btZ�Z%��`�)FpuQ�M�^����/�)���,r{�#�_���Ku�&�?"V��Tx�{4WG$Yw�H):R��M�4��p��s�n�O�T	���n��B��i�K����\0�bE��"���EՀ#n�iǸ��3Q�VE�"��6�>
��^4��A�vZ䯍�M�,*Lt�|3�F�Bڅ��%#��.)6��Z�-�d�v�U���u��頻�~��������3"�݅��K����"��¢HY�dr7��� q�O1����l�}�r���"���C�a�D��J��@��V�[��V���;[f�E���M�om*r��JX��󵵉�:_�T]�����{'�D���WF��X���w��Jt��ǔ��nd� �].B�����Hˤ�h]D�");�a�I�ɮ{�i���^�ޖ�W�F�����"��Z�eH���)b�>��n���a�>:V���6�>��zN �!SZM�b�>��� R�q��!�������q���.Έ
ʈTɯp��-'f���a����lwS��.��.A�����NQ�Elc"��F��.�z%�VFQ k�'UE�΋m���C0�B2�1�,�����.�N���+]���+>"v@���p���L�,)w�L�Vy��H��,ǥݱ��21�`D��+�D�M� z��.ψ*E�	N[���+q"�hD��E�Be��Z�'�4��k5�Ta�1ŉ.�+z�d�[T �5!jqW�)�P�|�)�M��qD��Jw��s׋���썐�RY!��«)�j=�dB.��bF��=���ֻ��wt���[���V��[Y�c#���t�9����n���	T�*tk�$e�Nq��mu�W�����<������\2�``&���67^=�M«˧U5A̷zJ�A3c�|m����N��2��4��H*d��PQ��G%�Zh/Gh��#ڦ�jè�������R) 	1��E{������m-��^m��L��Z�Hz&�Ilä� ��1��Cz��`�d�܎[�4RbtD�������bZ�!=�i�	�
��W��R$�AY�o��eC`��v�6�G"�>�u
":wi�'���v���@D����}Y	�^��N'���N�������-����
Y�
%Kz�XĪ5<	³�e�3[�af��3(�cv�Y�ٵ�e��0���aa��6��	�C�!�	։��bw�^�ec�Q���Ƞ���	L�p�.���y�[�OC���&��R�!�>6Lƨqj��`���	9�$�H(v	�p]�� h4l�OcE�f�ˮ�9��|Ov�����M7�MO��KDf�K�����/���	<7l��A�G�+&�/{)�7�_~��#_���yl�����L��6���2��
�},7�P,J�lA��1��4&�^�c�����AAlb ���aa���
v�P��޼�u����7�l۾iӦ��d }������_������G���H9��� ;I}ii �Ng�Q��$k���9+W�Kp�&�ѩ��!?77?���
uc%Π�9���m�扵{FaO�#6����n�:h�4q������P9�ʤ+Խ4ht�x敧8�\�3l����ͨ��3m��;�I�K/u��P��r\P̍��$��8�A�R�e>��U'2�2� �<�z�wF�)]}���d&�morȋ�������\���9�ڒ�[}��G�0};δ���}<�w穉k�J����~��;gHJ�Z�����}Q6���4�'X�ii��`dsY�'�,}�1>!�Z|g<�c�㓒e�$��]���$ϫ�d �Q)P���MvKw��EJ�P���6�@��R������,.��#%w�U�ȍOp�S;]F��xz~����z�,����:��z�������&SC��9���<w��ДJ3��z��U6I���@眚ɓk�.���=ǡl)�0�i �6�l L6�LT�����;�'����b��6���|U��<�6�s�^���o�XOd��6���:�v�����-cК�:��lw4ޤ5"�̇�
"�}y�蛖Gx���;b��Ӏq�q��Y��X�'�z��?r\��wB��[%,X>���x�br#k��Υ���:<>\�=L���C��Q��������,v��bW\�7�~��%�!�ɓ�E��:�w�*�5�j�*��cxu���g��|��?�_�UN����rU>�t5U>d�#hXԾݖ�,�]ʽ��ڑ���e1_�C�����A�\�Q�䒹���$ep,�n���8�ΜA�F[J�/�f2d���;R��D.�c8�P=L8!|�����.�
�;4�МGE8j���2��a��~�A�03���I�������ʢw��}���j�e�cז�k�x��+�{�����%��ݧf��,��D�k�'o��{�/�b?x��'.l=PVuD�#�: ��Š�S�׃��x�`�i�}:��m���cA�Y��1�{s3��@�<�g�+-�cg�����_���߾�����<���
/�%��RfB1�*�jUŰ�Iq���5���LZ��wA�&0--��3f��mO�R�Rk64�6E-f;��bp�3�foOx:�ҳ��/]�FNyt�'���}���KƩ؂u�)._��؆��<~��v�_�p�vG��je&��&�Q �ܡ�G�~��y�_`<�������w^M�9]��V?\U_�n�~��1o��_���Ԑg��8�x�u�G~
�"%�06��kփ�w��,&fYl$1{�(�)�<�5*�"Q[�g>�w�"��*��>��ݻ�}p�������Ҿk��lfvFy���ER#3��N�����T��U>��s���f�XSj6�|���c��-����LD>,o��#�X�ϛ�b-9HAKA.&BlC�D4E�J��[�QBRc6�9㘘8��g��?X���iT�=�c�����s���ͮ��S]ф�_��"d�����޸�:�rd��{b���r�%�Y�y;��S�<M~V~��l'�?���Ć���pϧq�UIw���E��_�Q��F�Ӹ�x�x��i������	!�]�jB�&U��Q��<�3zo��3W�L�P�e(���C<bw>
s���7��]ƾ!�O�g�O�������?��kي-[ZJWM`N�/ȫ�nO�����C��>���=s���=@e������$I	���l<���\��������������M ?#�I`U�$���T6��OrL�٬��*��`��<�l
u��E8j��Fᡣp�g�FW6Ae�*�}Ӡ�\��Ҽ>��v��'W����.����yòcS���߼�w'#��=�}��Tƨ��Q*�Es�aq��ڴ�${ߘ���=d�3"]3cd�,c��ڔ)B���lv�ٜ7�2{���D#F0b�@0�yY���dL�bOƷ9'Z{�d���y��4��Y����֦�?[��5�K1�ޱ~����?�	/i��G�-?l�_i�����t��W�����1�DnY�|m���D�g+z�{���|���5�>l 3��B>5o�;�����o�<�!Č��pl�8��s�a(�5���y���y�w��M������ױKn�����(!��4�0pРL�ΰ�J)��J��C����$�8��6Y��a��rڱ��p���:*;�b�ǥ�)v���V4XJ�#�k���xX.^P��U>5+X(�nr;4�6�(�R.��r�	#���1��'�٫�=)�/?�2���ۍ2_��)����d_�v	��CŒÁP�Ze5���86!�����Γ��`.���#k �Jn������t��ہb>T��MM�R�#6�ag����|n��	ܮ+G��	�G��֮*�}�B������[;��������ףz�"�?�iR�i�JpZ�Ƣxd��t���:�@ԘД��؄��Ֆ��.Q�KCb�(݆����8�hDP״~D�ITK3F�h'Nf�~��?�vZ܊��J?>�(a�n�����[����8���:���41~��`�/<��V<n�b�3}�|�# ZǠB)U�q<����u/���h�]���ոN�Ո���bƌ���+�#t�4;�`�@�L{?cL�}ܜ}�om�nnش��&TdPk��\<�Ed;å>�Bd0����n@j�̧S�� $ە�E��1 DLJ��"A_4�b�@�h�x��A��9�W/~vü*�ㄎ�,|��u��\�蕆*���!��ڊ��i�3���s?{�_�����FG��N�����IH4����1v52�|~��Q$���$ˌ��zh���J�2�����wLޱ8��	���Q�f��e~O�8�:��}��d�H�1J��)�i�i$V4;b�i�iy���7�?��B�	���mz�	~g�&?ʍ�p�5�a�T]���'pqg��*��ri��a!px��C �g4�0�c�|z�n����(
"@u��〒+g%�@�źX7�h�C�Ӷv�[�6����c��h+�`?~H^���:w8�cهoD��
�U
x��) ��$��D�3�AHxv���k����5�Q�d�F�E�IŲ�*kU2�^�Q�x��]��F~y�Ƨ'�?�̊���w�^�wk�ٝ�}�z��#z�B�Ǝ�Q���K4�Y9�xNQgM�&T��V�,4�K���vw?s,�mO�ً*��4$N�.0�-��r:ށ�oZ����֭��3'�����㥯�&����-���.W�˛�}S�%�6Ȓ�H�c�ڴ:���i�*c��S�	M<��DS]��6$�b<�>�q=�a��g�I7V^rw�9yeGvW�0� �*�!-�& a�Ѳ����4��B���� l�ږ��96���NL2l�O�g��<؝�m�Am�����ST���S�B؛	v7DJ2�@Q���}d4�� d�@����co"|��EeAI��L|n��ZZ����w�^�(��������fd�����M���cĮV�%&5Y1�����&k���Uа�����Vk\�	5qN�2�F�����D�Ō�G8U�qW�	u�%ځ��q�37~{9餩e��O<���c����N�$c�{`�az�۟~vn�<}�o|X�7K�V�Tɢc ��p�#�-=�^Q�����q����9�۳cY����r�xVa:���!N�f���S��*w�
?���:�%g^z&u�/����7�\�>��)�=���PL����AcaYN��:���D6Z�-A�	�5�g-��f��QS�눣���>m�'���!��Ou�}C~��	���o�����C�:�۸���x�/z��'�&t�̞� h!g��g����,9"�:؉�4z���ӳ��f2�g ��1zk��e�I%�HD��^��?9��k�vҀ{8w^n���R�I�/=�������W�܄������N*��1	����ș�O�U�5�1�g�d�_�1�R�*���{��@���G
DJHĳ���s��`��Ȗ�;���v��YН�[;r��&�C����m��\�f�AZ;�t����Y��47p����T�>�}����*�M��z큕O�~x��L_�K����z��=��7��w;�^<��g�?���n��`���z�FéUj ���!x(�g*֭*��*f��;T~��u���:��v�.��e\-?�Z���)��(L��'�5<�c���>#�!�����e.	�A��.��K�#{�F>=��(��c��D�w=�o�h��.�}}��%9xn`V_}</V����XM�O�F��T�jO��]9����8� ��b{Į�ݖ��&s\�����qG�"O�|~��G
�Y3y��_||1�Xܦ��/.Z���07����R��_�쭼�mPP�8n��#���'#J�w��ɍ��Λ����w>��K�F��}������D���WWG�:�=#��s=q�jU>�Zo
w�ˀe5��Xxgz�������G�'�u��O�g�w����ff�|@ތ��T<	������w\���/C����"�4�?bM�Nk�Bē��n�.�ǘ��b�|qq�ZS�������dwi���H��"D%_4�'���Ps���O��k���e�yW>�%�/<���8<�+�믷�v|6@�e��^[�b�\f��kNN "���K�%�|U6�l&�em6V�1�|F=6�z�Fźn����jkg�B�;�a���3vzV�":l����e�����}y���t0t�oG���p�3-ۊ�,c���K�8����9�����v�YX��/Qڷ��,�M��� �b������G����7�x$������x_���
� ����$ɮ�3_b�ݚ���n_��1^�U?C���`H�4��&ead1X�ׁaUq�jU�*1�5t��xȀ��|�#:Fǃ#�q�M����ͽ����>6���F�^��b2�J���(�?��8,�����J��zs�����?�Y�������k~I��07yZս�LŻཇ�AIr��p����<�Rs�=Ұ�՜EA{> Ip���	|bAN5$5p�?S�ǟ������Vy�9|^�-dp�Ҏ|fd�[̛���L�?�#'�j�F���"������1*-�95od��y��{�D�y,�c��O�o��;���p&pZ���1���d�t�|Ǎ�������@n�3IF�NǱ`�U�q��q^��&L�Xw*9�3�=y��Ͻu��^�"_�/_ƯC�i�G�_��н���J@����~���'9Y%���G,TFf��l1�v��(�u���r�������ڤb��:��]Ǡ�ߎ ��t)`O��y��/m��Em8��y���N�ɘ+���;Q�k��q���;�u���8���������Ǘ�^��n~��c�Z\2{�a���Y�$h���F�8�A�i�t~MuZ-��*�Mٟ�)��b61i�����ɓo����'�������\�'~�`=~���RJӱ /+iL�'%pjFê�V�R�Zr�*	D{{�a]*��a�b���;lnG,{����#��c����oX�I�0��D��"� ��a�t��w����,u�0�:d���)n*�X|�$r���Rc�q�/�e+H{��X;{�@�Ff{zf��<l�`{�����4��sx�S���cۨ��Jn*{���JwsXk�5��g��Fn'w��XN�8�������2\��0W��b���T�h��� ��>�l���2ڼ9��n�q���ڣ�3k}��(������>I@<#�y���i���4��Om�P��)y�9��g��<ÏG)h�͑�QgƤZ�%&%Y����ج���~�Ȣ\���:o��Y#�������jx���$��u�M�!�ƚ]����F��c{:-�E!��y�i��f�*��Ē�~q��84v��xŗ�]�����>��Č�/<~`Ⓡ~�2�����)9���R_p�3��{u���E҃z��k�=��[Gl+Z�{�%�%}��3.>�cZ���z'͚��\�_r����Z=�ҟ������˪�#�c���W�;fɋ]���)O�~������<aOǶ?��w��s��2<J���B-p@��m��#�t�K�zԌ6A}6z��ы�lEG����6@�(*B�a�R�w�
�!#9���j�Xo�:��f������\�Ƃ�	�O������?xne8��Y�D�l�����嚹}����	3�]��*�j�������Oi�L�L�1����z��u]_���3zA_�ߠ?�3*�%揆Q��yc�q���ę��L���M?����Bc���Ѧ	e��@D��f�Sқ���xo7M12B+�T(��Y���*e�<��y��T���U�*��)e5��]��5� j-k!���u(�9��_Y�y���X�R6�6�`�i����)e��!���d��J�E��AJ��1�̣$n�R��S)���u��F����AI��������V)��]������>�Y)Ǡ9�yJـk�T�0�!ܰ$P+���~�&ش��av}XL��/����	g��c��M�f�!ؘ�s�\q2,Q�g�ck�Jf�c���������s�ͣC5���@�8P�c��{�!R��������chCH��fm`���Wb��7bs`vC(h�ƆF�"�<K,��a��X+N�8����&@k�a?���9�B�5Z(���(���p8
6�C 0�jhd��j�Ņ��X5�n��Y��޳D���n�`�0�9P��74�C�Ɛ
47�)K��z��}^ ��P�;w1�m^L�|Z��'� �	��{����aņyM��с���@���k���6�a�z����k�	Q� 5�&�������  ;�����(IC��!:�1����V��$ <7��R]�Ь��w]�1S������̟G��w!�iB_�\V�ʪ���gg/\�0˯�ؓ+g�R_xqS@aI3Ye��R��F¿���d�cKŉM@/ '*2�.��5Hdlh
��Bs��ͳ�'zKQ!j S� ��N �"n?��P�ބ��'��UD���޹(�t��QA��E0�A�D�~�n5�,pc����Bi��E1��	��0�V(�y����"O�A:o68���یF��	@O-�!��p��
��{/�	u��F9��B����˫6�J"�q��,�Q�mAp��D	�(�B���Z�*Y�F��Qet&�B�Bk����ĉ ���Pv���kY���r�B�9@�f�A-�׵�@�w���T�S�P��i;��h_�Cʾ�4#ķh�vB����]O�~J�Z���Fe�,�9�a��\�Fʹ
�h��u��p�e?ݵH�%���R�Oy��<�ӱ5�>>�m�4�B����B�����'��4� ��ӽi��:Eb	T�n3��m��\"�	P,I�O�̘K�F�r�\(\S컨V���n�-i�Lu>�Pv*؊ҟ]1J��RJ83���v#Ŷ���)MF�U Ew<�ڤ_us��J^���t�����u�6aj�bT�(ߣ���)�����Q�O�T�5Q�Vp�G5���a�e6`G>YT{�O��=Y
�����^M��=����y�c�b��o~M��D9X�Rj9���*��X��Ν�s�t�.��� �0�'Di�E�0�'��h,M/���g�ѩ����OV���)Ȇ���NxOD�v*p)�I�H4���?�wC������-N4:F&�zgA��\0�-��pG[��h5��m͆Vx#��pCO��48� F�x����yu:�F�q!,@�Q��X� �J=꣤��W���ƛ���w��7Ϲ��Ϋ���k�1'��]װ�Zյ�5]�.3�K�N�_�Lu~��H�W_&;�_�>_|�u?���^��/��?�x�"+]��^��9�a�- �*�G�F��ⳑ�+�hv F����ö�n��W��R9���3>_!�/;�r>r�3���=Ϊ��o-{�=q
�Y��l:���9�Og���g�ǜǘ�c�ǂ��p�?�?�)�紗�7������פvk����i99µ�f���];Ķ�)co��%�)�D"'#F����]�#����?��d�����|����^ft6�\l�} x���fa&Ɏ�vT�h��nے���7ՙ�U�� ��8���������]�5��F'�Gy{q��^�|2��i�|`�ͬ��� ��ّ��k|"���'�=q�	��֣ �K"���T�c���p�&�ܔ��	nZ��AMō,��yc\�Wܐ�����j}p=���9�e�c�u&��t�r���ΓXw0V�%��d�]��\3n�s����U�p>:�ӹ�lzX|8�a6g%^�K+4zo��j�;�U�{�*T�B �VC_�G;/b�Ag��$�5�;sZ��>� �txO��5�R�c���eA�ՇG8�,>��q��<����to;�J)���D�I��iR�]^iRJ���2|��z�8K��βv�(���c�b����_�^�2-^���\{�+L��
4�~%%�:��|c�q��3���A�F�c�Q�m׌l�������xS۔򌌒vU�䒈�lz������4iZDXAӦW�a��������OI$��2R��W���D
-P0�is�_(
�ψ^X)�PFF8oZ�=p����
���!�f@-�1�>3B���d,���C`MaR8#���f�0���GHXif(���L�+���t�63�4��^q�oK�U*
endstream
endobj
xref
0 14
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000392 00000 n
0000000115 00000 n
0000000549 00000 n
0000000604 00000 n
0000000761 00000 n
0000001869 00000 n
0000001901 00000 n
0000002622 00000 n
0000003053 00000 n
0000003253 00000 n
0000003833 00000 n
trailer
<<
/Size 14
/Root 1 0 R
/Info 4 0 R
/ID [<536835330C477215CD49D6A1AFE97232> <536835330C477215CD49D6A1AFE97232>]
>>
startxref
15263
%%EOF
