%PDF-1.5
%����
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/OpenAction [3 0 R /XYZ null null 0]
/Lang (en-US)
>>
endobj
4 0 obj
<<
/Creator <FEFF005700720069007400650072>
/Producer <FEFF004C0069006200720065004F0066006600690063006500200036002E0032>
/CreationDate (D:20220919020032Z')
>>
endobj
2 0 obj
<<
/Type /Pages
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Kids [3 0 R]
/Count 1
>>
endobj
3 0 obj
<<
/Type /Page
/Parent 2 0 R
/Resources 5 0 R
/MediaBox [0 0 612 792]
/Group <<
/S /Transparency
/CS /DeviceRGB
/I true
>>
/Contents 6 0 R
>>
endobj
5 0 obj
<<
/Font 7 0 R
/ProcSet [/PDF /Text]
>>
endobj
6 0 obj
<<
/Length 885
/Filter /FlateDecode
>>
stream
x��Wˎ�8��W���ÇdI�b�������n�`s��O��t�jy&��<�*�E�$S�ݿ�:�'���ܗ�]*��o�>��no`|�|/�8��K2����ս_�c�.�� ��ǟ�/��r�P�c?TBR
i�D�
�I�0z�X>ь낱E��e�� VXML�
��>��r���	�%N>��̅\3�{#OMӉ����3��0� ��a�1�Z��(�*��H���s��ʫs,�B�	�$��$�JB��(I�ˠ����V� � fq8Dd>Jv@%�	h��vw6��@���}x�B��j��xGR��(��3Є��fx3����J=�梡N�e�F)�� �VC���jeB��k�b~+����i,�^�����K֒���|���׷3(R���|�B
9?�*g1��6.��
��Pj��(�b9X~ Ȥ,�YEU�F̫�@8���2���fb��&o��05�D�bځ�f߬&�=Di(ل��^
K��C�M�>�'tvw���k�9}3b�{�|�^�$@0�� _��Gˡ��Zin��\S�}�xф�h�qKϖ�W&�J]����*6-H�q��q�,-���\�D��@zv��Y^���t��-S>{�ٶ�<���1j$b�	Xyj�)ֈ�e�H&젷�_�����L^H|`(���-��yr^�۵���w�y�y�Z��h⏹����P[�U�n���Y��`���&�4�측�`����~ī�`���MJ�iEy5u`���%�?)��T������V��/o?!���e�r �8�ך@dw@����Bv^?$Vg]�����Fb%}������w�������9@_v���\��=�>{x�v_u;�nɯ���C�bF
endstream
endobj
7 0 obj
<<
/F1 8 0 R
>>
endobj
8 0 obj
<<
/Type /Font
/Subtype /TrueType
/BaseFont /BAAAAA+LiberationMono
/FirstChar 0
/LastChar 62
/Widths [600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600 600 600 600 600 600 600 600
600 600 600]
/FontDescriptor 9 0 R
/ToUnicode 10 0 R
>>
endobj
9 0 obj
<<
/Type /FontDescriptor
/FontName /BAAAAA+LiberationMono
/Flags 5
/FontBBox [-481 -300 741 980]
/ItalicAngle 0
/Ascent 832
/Descent -300
/CapHeight 980
/StemV 80
/FontFile2 11 0 R
>>
endobj
10 0 obj
<<
/Length 490
/Filter /FlateDecode
>>
stream
x�]�͎�0��y
/��Qb���H��Ab������H%�LX�����m�.�>'�ן�����;�ÒSw�9c�m��Λ��cf��nI+}v�v�����-�z��j������i�O'�)˿�އa����c\����_���"[�M�ϱ��v��^}���}�<,���_��c����R��z��·v��lUk���י���Վ[N��gb���E�v�Ȏ\�E�p�\��Y�k�F�����;��5����l�o�_���o�;�ֿ��f�>.�-�%���2�>���>�����OK�-�E��_p���h��O����Kdb��hO����ҿF����ѿނ�_���?|\��L�Fk�_�.�l]�����K�J�ҿ���w�t�/�&�5�/���_����p�пBΒ�q/����_"CI��,��L����$�]��(��)'u����0������5��C�c�����F�w��i�.�� ���
endstream
endobj
11 0 obj
<<
/Length 10865
/Filter /FlateDecode
/Length1 16348
>>
stream
x�պy|U�7~om����,��4Y {��	�IH��I�%M�!aB:�; �Pª���"* He����Fg����m�QtTH�=�������>�?ow��.u�9�{�=���	����!	5�����!��E�j����&��Q/�5/\�䱹�b�"�xya㲺ߥ��B�"��L}�_���e� ��а�� �6��_�'�tF��Pok��]��@(k�/���b�P'�|�q�?�u8��DH��9
�D)"Bc���h���j���.�6_��B�#u�fXN�T�5���`4�-V[l\|�=qP��wvINIM:,=#3+;'7�=<��Q���1v�x����=˞E���Ȋ����3Y�R�z.�Zϥ��hY�%���)�2�x�����m(���֡�ѳ�k����ڈN�h��:+��6T����}(��A{��@�U4�cU�0Z�:����`���E|��U�^�N=2<�>a�����>���_���w���55Q���h=̰�*��7��T��A�a�5�J�h�Г�Zt/�Z����ov M�u�x=��4���4C�>B�*A�h��EtTj��;��O7S'(e��a�N�o-�ū�.�O�w������=G��bj
��\a}�[Ԅ���A��h��E��I=�P7���!��К��� C�`��{z���b9��gl����Uq��zda~/Y�ĕ0�O�.^ܐp�پʊ��3�{�M�RV:yRɝ�⢉�������1f���#�ss��23�RS���;q�A��ѨUJ�24�Q���:�7z��b��$3�/��/��(vy�#�����Iq��HM.���#)���k���f�mo
�7��7����.>r���w���+������#����̤H��8�0B��H�G<K�ۋ�AFܡQOtM�33P�ZE�"i���6K*�xL��1�-̴�_�N�,.�;��̌I��H�B%�nbD!����hߑ�վ�ӀT�kk]�����c������czd��(2t��q0�@$�UTI'TKg��)��G�d��o��t\�/l��-\��;D�jbϨt���X��{\�������Ӷ��\�Zm{s1����@�����g�/b���c|��=3J#��s*#T����C�����Nc�;��ԍ  v:	:� *����:�؏ !;���IOWo���������v�nK�+�#L�ZW1 ��i[ ֵ�(�e�辷;]�&#?:�'�˃T�j�� ����nȐv�T�}}\�����2�N���Z�[Rx �$=j3+#B���⎜l��5Iʌd��#Wa�v�X���yX�21��k�Q��bi]����EQ-������s�c8o���WD^�M+K)n����8�����J�3"�@�>We�G�z�.�O��������+GɂD;9&��62�J{�`D���+);���{��*��"Y	� �Z����+���bD��Ł"�=R@�%�4���G�@gb���sF?�t�2c�$���v���%�����`G���t\>W=��dn	e	sYW3���0!'t�V�O��?��;�z_���I��|��UZ�N��d�$�AĄ�QF��Ȃv��������!d1׏!D\�j�]�c�����g_Nx�P).�Y�����Å�M���ٕ��Yy�����B_��<�æ!�R��4�
O*���(����2�^Fj��5�Im��6�j:�h�!�(Eb$ 
z�h���6m�h[��&}:�LP��RP	Z*��w`�tZ^�U��KZ��0j��܉�:T�=�F�!D%\Wq�u��ʗ��Iw`TH>`.q��l�V��Zb(+|���>�ؐT8�]�AM�� ���]��UH�H{A��#�
0Ql�0�t�`bs*��$��3�v�e�)8�v�W� �J��WQW �P�$A�!�h��%Ax���sF=��6�ss�F��v�+ij�C�+�&j�h!���ߧ栗�N��E�c�/c���KDrsp�ӊ�R9��ݻI�w�%f	;�P@(0�B����8�3�(�ʡ�bX���g4���pG#����"���ii�S��*�ʌ
ҍ��]5����t�y���m�K� 6��y#F�RNNެ�®��B$�w����#��WT._�/�7_x��/^��x��/��T��1��D2�� �$f*ҠX�&XL�q(.^���T����6	���C(�g$b���)����b��I7.��_��~��O�غu��T�>��`����?į������O�H���Z��������T0J�#I�T��TiC]����lz�A�w� s(��+(p���>i�k����q��]���X�{<v��b��5�M�s'��s�q�������TZ�bIݾ�	�S����ko��t�k�V��ͫ�]4���٤}߾�Mj���YL!��\h�0(��!�l�{}F+ȫ�SN��� <7A�N�'���sp��&�DE�g�x��,s�;����q�[�_Y����zl�rjp�;�ʧDK��k�� �/>���>~���6��:�w0�F�L}|�I����	z:'ה6�g2i������W�{�Y��h��Z��Ǣ�>�Uj�$��V '��Mf+����休V�58%ե�L�7$�̗�H59�
,���xV�(�"3%�Ytg���б�����K��K��'�������m3N.YQ�*���|�c�;ͬ4�!�v�Y����'g �953fԒ���T<�9e�D1(Nɶ�bc��f��TPp��n=IT�{�d6tmChŮ����St�?���{���M�F،��νz�;x�]��2�тݤ�Q:���Q��V�N�bj=b�>d�.(0��[�ȃ����|�����;�:��L�Kɚ�!�$���9��x�Iq��8K��[�*����BRm���œD���>Y�?L��B��R�̎9��s�-�-kٯ8A.|��ŋ8]��֓;�h� �w�%�`U*D��
DkcXe���f��nl��=̞g�e��2U>�tUU>d��#htԿݲ�-[���ޝF�쮥1[�S�����)��h�X�$1��	6=]Hgh:�88V�r9�v�%�답t^�ZgE
��gr�a�y��	�}�>�ݽ�lwd�Cc�d�Q.d���n0g��'yi<��;��i�{�T���u�ͳw?�I+�����?�~���_��#V���/���8�p�a[�cM�?i�vā�o}����>u~�ao�1y��u �[�Ac�F����aY�^�.�i����#�����Q0P���h�����|���;^qs~N|��ۛ7o��6���|�֍%�iBFB1�"�lV����8���ũ�5����rT�9NM�C��y�t�_���7{Q�ъ�+8)\��ƅ;�ʸ��%�ǋ����R%��_�}�7%sŃ8��;����q���O�b�� "V�׊�
[���3��>�A�� ���8�ѷ�SR�d_��y������^�ǿ��d�����7��P���[���ܐo�q�ɞk��L�9B���,�-֨�oSB?xLL�XO 1�e���%��ns��	"Q_�o<y`�=8"z+�=���={胛q���������o�vEu�G��b�DF�W�&3S� ���1��۫�Pl�H�6��c#`��s��f<O��>��l�G�R񨸃-��/c�?o|��� � �����h����5E���A�8��s�Q1q�>�OYa��U*}ȧR�֐���}�'��u�횤p�7�p���/�H�e����ׯ��/۴繇ݽk�Xy�zF|Q܁k�L<���Ã1݃�O�/����6��R\�BU�(�2icc�I��!�V�w�w���{�����i�5!�*hU�׬hSP
��;{��i��e���7�j)z��n��v>3��ן�]���O��N�_�����?��{���o+[;�:%>'�ݰ�����^�z�}�/�y�̋�.�W����|�-�H0M����A��z,�-t����Y�?�Q�����GG��-��XKS�ޠ�B>���G�C>�<e�B�}ɥ��:ip'���2��o�d��C۰b�s��0�=5�mu͍��%~$�(���%�!`6���\�!�~�3RMF�1�Ӄ��M&�9h��	�;%��VEn�t����T!)��"�� "$!��
Jq�����q>�CoL�-���қ���ž2��혳�_��-3�<��Q�Q˿Nt��ۏ�WΞ>a���e�G�]碥˃�C�_}~i$�1�9o���sJ /�KTXt�AI11F�:�3*pJ�q�lzg �<��IuX�n�}�Ȯ��m-�b:-WN|�������к�ϛW���羻�~�	}u���駋b4U
��qf��bQ*bl$]rX�C>��n7�|v;c�����V�d$�8w"n� y��"E}�!K�2���I Ŕ.�b�}��v��M���0���H6��^3��ų7���>c�`��+��I�������[(�<5�!U��p�REA\�u�j��k�lmP��N��8�J�ռ��Bl�R�����lUa'������ߝ��Z|��X��^~s�fzbw)��)�!dP��JѴB�%Rk�B� �E���kHB|��e0�a�e2���}��0�tWv_�
ʏa�Pda2g���W.�P4�A��=��u
Li�*�V���ĥJ���ٓh*��yD޲ p�r��Ur�N�I��[��J������7��?��������C�~q5[�ӫ��ԏD���@.b/q�D���S*̆���G'�3�����%hu��Ri��:Y$Ii�� ���)h��j�Ͷ�"������ϙ�2�/�f'd�]�����
q2�m�w�n)6����?���y��!����0�0�ބ⑙cR�Zm�vBs��lZ�%^��k��>�1��)�!� ��:$o���i�;w�$���w���s����X�  ����3��h�Y�]�ܥ�l���<�j��i/��'L�?�ܚ�����ǖ�iS[Q_l=��AEB��aX��hY-�{1^�qƘ�P�V%�@�	I��W@nra�3��J7���-���p�3�`:�,:8��6���歫�j�"��{�f�a?�A�8F�B:��ӻ���:��>��@' �to.Mh���iʱ��˩�l�uh��/����{��s�[�L.E��d��,}葍k[{ϋU�Q#�Z�?sü�>��?����ӛ�F�A��g�{�:�J��V�����>��ƨ�PTorjċܿ��rb7��eG�e�t�ع,��
�<���u��>�~p���\�2@f�X%���ԔTcm������|z"�7�=�F����8�:z���G�͌œ�3v�g�ͬ���9������Zs	6�5E��'���Ð�&hc��D�?TFݙS6P+1P��V��e�'̽����%ˮ_��/�o΄�2����ì6�~�z��l�lЊ��WH��u�	�aC�A���5�sB��l�L�$E�����m��f��qA"�C�H�x���f�	�3�&^�.�������l�~�/8c���M�>�,^��۰��/�o:�����Z\�r�8x���q��~�#�2��lQk,�͢�*�^�0 $�G�w�)x�}>���U����J�?{V\~G�9�����xϵ`�j4\H ��Q*5M�)�FE�+8\�":#봠�/�u�O�L�|������Z�pW*���;[�P��b�*)�6NZd�\)�� :`9�R_�SҜIڂ�ү~�Ove'��<F1�	~�Z��ſ��g�`�K��^|���7��E����b��G�Vq]� �B����V��X�3!��냐YI�|�10� �٨'͏�@9��.�7mo������T��o'��a�q������H�t.9
�T/$� ���d�'6�12���fs���̩hi��I%fs\�Uq��J�� �o����[�czխDD��l@}.^>�����S�{)��ж�G�M�f�ɘ�o.��QIX�ަ����'��[�X[����2yM)P�`R`�P��MV6�.e+�_'�bf8���,f�Ν����8(O��e���-�B}�f���$c˓��;b$Xۙ�D�,8��2��3l���w���j�!�֞�}@���bbTX��u*M3*&֦�L�L3a���4�2]5�Z���%����Ʀ[�m�ވMJQ-���� ���ȕS��_�7x����5��	���u����;���}�8����Kg\8�W������=؊b=��פ�,�V3N��ʄlL��j9���i�
�zX�ALki,X��`�*�ʧ������r눃h�d�0+^E��{����/�����-�)��-�:�"'ɼY��4�e����CR[i����b��T���e��x\��׮Ϧԋ��3�[���{xl݃��.��_�_w��kG�g.��	s��>{��'�}��Q[}����-$r`�
p�*�6�Q*� ��� MD�Ӗ>ӕ�|�G��ޡG�o�7��⛀Íow�db�s\->F���!��O���)U,�s���1#�`COOO�:	ڠR��Q\���3�S�Q�w/��2�,M�8v�mP��D�df����|�oРx�VU���QG���|w��	OK��$��R��~1!o�$Q�IS/~��8r���ȣ����hM���g����.d���z��U��e��W���wq]��-��Q.��ɇ^�q6>[�˛\�cg4�|zn�a>�y�
*�E�W}��9�DS��`�?~Z]��e�e�EA�%+ѷ�`eHə+��/��vCT8k'�j`W'��X��A:�ŪtU>C��|��9c/i$������N��?B�t�+ψ�o?��3ۨ��aq�ó�t0�g�������x	�6��{9s��8Dk7��U�I�+;{�	�1ƒ��*_\�T�T�4%CADBɒ�
�����{x�$sQAɏfd合u�H�t�)_��'�A�Uxv������E�d����k��!<��w�GG������φ�ػ�����gLs�<cR�Z,�6$�y~�#��B�i��V�t!�^���V�R��['d�r�o� x_JB���SV�L@Aֿ���ۏ.�Xy����GB];���,}�����ɏD����\�B�����s�.��u�ĥ��>�O�~3̇�H#J�*N1�
���R��3U����{�lfܗ7�r��ɧW������"��⛇�����!<�`��R,?[��Ȥ���C+�╊x�=���4��x�:�&M�f��Ұ��I�lqF7yJG@�B����N#�.:��n��:b��$���SP�:�et��;2ϙj^��j>V	�\ ���Ά�@�������#�>qVCc�쪻�*	�! �~�G
��搊a 7�]X�2
%���"�1Xɘ԰�
@H"Ӏ�x�v�")�K�sSux�9q
����.n8�?����(ܽ������:���>�_�iȯJ�J��C#ǲMk�1
5�%����q�c��,ѭ7�V�������N�]b�w8;#��^|B,�2(�8?�}��C����཰���%��C��V��j����~?�L��r�;�Ɍ�@�ɮ���q�� e/�E�.�W!�3�c�.���ݽ@����F��؁�O�}
vA��@��m&��ٮ�7��{��=�E��x���p����yM,���'�Y�0�;�A�8�#���.ȭ�hN0YK8ZOa
e�#�"hl\������U��a����ѳ�;��=O���?!��a\�̢/I��]�V -��a��L����b3l�&[	8�C���ո3^���~C�'���t�)��(."� ��r�6m���D��?�$U��~G9����������_d�q������q���'��k%��_-1s��S�t7Z�j�K��B����-�]��A'��mB-h�n�k!97C����ӎ�C����9�A�@�b�=@�4�zWî}v�:�m��㻰4G��!h<|w���#p;�P��:*B]�����L��d�l�}�}�+�r�Y���}����;��Ty����*Q=Jݨ>���f��Y�G�֤��ݭ�c��P�ޘ�ucu{u���[����PhX-!R�r`��c@�h.���i#h��&�>����#=԰<J�r����Q.3��Cr�E:��\���\V��C.+�b�hY�t�@.�a��"�5(����O�,�S���i�\֡��HϨ�v���e�� ���)�c\r�FÙ\���;�̢D���Ay�\V��̫rY����rY��?�e5�5��\֠Q����Z4We��1h�j�\֡�?5,l7,������	6/kiXX��j��y9�9������ ?1��l��MYꉷ���� %�p?��&��aA �.?%��X���o��	4�Z�L��n��h	�r^VNN��V�m�6�x?n���[~��
��6�hlh�+�ʳx�?h
���Z~f��iuu5��&�����p=ȹ���!T�PC������Ey8�$�O�ÁP���^ ��`k��)��/�o����C|m ԰�	�,�����ij
.�K`XK��%�ohZȇ�M!>hi��I��z��}q ��P�ol\j[�C���6��	���tj`遬^i �: �oX��\"	��i	����ֿ���!���-���k�	I� |��)���%� ag�Yv�E/
i(ظ$��n
jCD%�0�F���_�)�[@��p}f?��Ma����0w ,XӺ�(��
�i	B_s�?T������1��K�.������d��_�/k�*i!T7��4��JJ&�(�T�Ok|< /�����gnV��`lh��B�Y�����<e�5��n �� '�j��~(ՠ jF��œ�ꡕGi�:�y�s��ѝ�V�a<�&B�F��_�DM(\���OjyP�!KQ"�΀�$_�`���O�GS�gP���F�mAP���V��L�~��/��%�����@��f!�ώ�e�@��0K=D�Œ係� l����$���' �j%��v�Q.��F��&魙?�qp���5�{߬�h[�RB�^�s`�"IP+��[8�;�?o�tK$�S�vRI}�P��bFh�Jh�v��R����~	�Z���&y��9�y��X���&IsKdI����u�=$�m<��ҬyIZ�H�mR�j~IQ�/�ް�n�7�w���FQ����TZ��}�'���N��R�`I���ZP�l��+��"�������|����V��(��U/ى_�r@�zX���Zy��w�Ԓ	a_�ĳY�K8�_Q������R��FI�P?�M���R[�i�V��):�F�'��OKu��EѬ��e���$l�2נ$Q-|�z�ZXƶJZ����]��9��oP�,���,�bi��Kv،�@x�ґo�d���O��z�d����#r5K�_%-}�,�d?�Է�Z���^M��7*�<G�l?9�6
d���=s�_�m��Zc�Ò<!	�,i�p(����Gt�+��τ\��T�g�ϻ�LdA\O<�!7d7������s,�?�w@�<���#m4!G�(�ʂ7*�y�j���኶�¸h���m͆Vx"��pA�w^*�p��*:q�q���q4O0�" @��@`"(�g�\/��xaa���y��x���s\��;�\�u��:xu�U��U��*v\���J�K�%J}�����)�������$��K<��=��X��cs���q��{�_�����8�	lA�	���8����?W|6��
4��m ��0��p�0-+��E!�&�F���q�Z������ȧ��S����z#���7�S����G�I̟�9�u�n>�v�ҟp���O��8|��	���ߙ���l�l�d�/@����1��k;9ƴ���/�t�%���Jm��*銼���v������>Xp����:��jB֣<��y ����a���;�w6蘭x<��kO�#g���^zܖ�!���=Oo��=A���X��;�i����=����Nm��m�r=�6�nZ�G�h����|�꣬��EA�x�M)���{�✭ر5{+ܺr+����[h�'�-q�~s�fjڦ�M�Mt�F���ؘ��6��)H�y�r�{���H,�9N
��`�lX��X?y�c��q���u<4�Ǳk6<�?�� �� ^��UZO��j�+�UĻ�*n���VC_\�{.`�G�G*s�g���\O�c<g�Ӝg�`1]���`�ʣ��=���xw$�!t�#6�Ӊ�B2��;�N�N	��Gy���i����|.�r�zJ�Nl�ɠ�I X	\w�u؃�{�z�6���
[����<}+��J��:�}�~�������A��y}�^Q mW�t����m�ŝxk������NEό҈�;'��E���]�>;­����s*;0��[�i*T�+��T�Fj� �B�:l��
�­����!���S�H=p���&�
�Cr��Z8�U���B�ɻP@�ȇ�� pz�>E��hFҰ�zY���t4?$U������'��PT�P/G����t>Ȁ
endstream
endobj
xref
0 12
0000000000 65535 f
0000000015 00000 n
0000000288 00000 n
0000000386 00000 n
0000000115 00000 n
0000000543 00000 n
0000000598 00000 n
0000001557 00000 n
0000001588 00000 n
0000002001 00000 n
0000002200 00000 n
0000002765 00000 n
trailer
<<
/Size 12
/Root 1 0 R
/Info 4 0 R
/ID [<92CA4A2A10B36E88F4695584F96318C3> <92CA4A2A10B36E88F4695584F96318C3>]
>>
startxref
13722
%%EOF
